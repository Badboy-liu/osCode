conectix             ;� vpc   Wi2k    @      @  �?   ���raWo��ރP�ϓ$�                                                                                                                                                                                                                                                                                                                                                                                                                                            cxsparse��������             �    ���}                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        �      ������������������������������������������������������������������������������������������������������������������� ��� ������������������������������������������������ �������������� ����������������������������������������������������� ���� ����  �������  ���������������������� �������������������������������������������������� ������� �������������������������������� �������������������� �������� ���������������������                                              �3��м |��PP��� � ��  ����<�t�< u����u����L�����t�< t����< tV� ��^����� � |�W�_s3��Ou��Ӿ���}�=U�uǋ�� |  Invalid partition table Error loading operating system Missing operating system                                                                                                                                                                                                                                    � ��?   a�                                                 U�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                �<�MSDOS5.0     �� ?  ?   a� � )�<NO NAME    FAT16   �3��м |�x 6�7VS�>|� ���E��|�M��G�>|��ry3�9|t�|� |�|�&||||�� �P|�R|�I|�K|�  �&|�|�H��I|�K| � �R|�P|� r�� r��� ��}�u
� � �t��}�_ 3��^��D�XXX��GHH�|2���I|K|� � PRQ�: rذ�T YZXr� �� |��.|�$|�I|�K|�  p �
�t)�� ���;|s�6|�O|3��6|�%|�M|���ô�M|���
6O|�ʆ�$|�6%|��
Non-System disk or disk error
Replace and press any key when ready
 IO      SYSMSDOS   SYS  U�����    �� 	 
  ��      ��        �� �� ��! ��# ��% & ' ( ) * + , - . / 0 1 2 ��4 5 6 ��8 ��: ; < ��> ? @ ��B C D E F G H I J K L M N O P Q R S T U V W X ��Z [ \ ��^ _ ��a b ������f g h ��������m n ��p q r s t u v w ������{ ������ � � � ��� ��� � � � � � � � � � � � � � � ��� ��� � ��� � � � � � � � � � � � � � � ������� � � ��� � � � � ��� � � � ��� � ��� � � � � � ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      ����    �� 	 
  ��      ��        �� �� ��! ��# ��% & ' ( ) * + , - . / 0 1 2 ��4 5 6 ��8 ��: ; < ��> ? @ ��B C D E F G H I J K L M N O P Q R S T U V W X ��Z [ \ ��^ _ ��a b ������f g h ��������m n ��p q r s t u v w ������{ ������ � � � ��� ��� � � � � � � � � � � � � � � ��� ��� � ��� � � � � � � � � � � � � � � ������� � � ��� � � � � ��� � � � ��� � ��� � � � � � ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      IO      SYS'          �2� F�  MSDOS   SYS'          �2� ��  COMMAND COM           �2� u�  DRVSPACEBIN'          �2� � SYS     COM           �2� �$  ATTRIB  EXE           �2� �+  CHKDSK  EXE           �2�  �/  DELTREE EXE           �2�" g+  EMM386  EXE           �2�$ ^� FDISK   EXE           �2�3 �r  LABEL   EXE           �2�7 �$  MEM     EXE           �2�9 �~  MSCDEX  EXE           �2�= c  QBASIC  EXE           �2�A � UNDELETEEXE           �2�Y 0g  CD2     SYS           �u!] x@  EDIT    HLP           �2�` �E  UNDELETEINI           �<Wc �   C       BAT           uQ�$d "   HIMEM   SYS           �2�e �q  CONFIG  SYS           �b�&i y  AUTOEXECBAT           ���&j -   MOUSE   @@@           c��"k    CD3     SYS           a!l N  EDIT    EXE             Qo  EDIT    INI           -�lx �   DOSKEY  COM           �2�y �  UNFORMATCOM           �2�z �1  TREE    COM           �2�| !  FIND    EXE           �2�} r  RESTORE EXE           �2�~ ƕ  SETVER  EXE           �2�� �.  SCANDISKEXE           �2�� f� SHARE   EXE           �2�� �*  XCOPY   EXE           �2�� "B  QBASIC  HLP           �2�� A� MOUSE   INI           T�"�    SCANDISKINI           �2��   MOUSE   SYS            �� �{  CD4     SYS            ��$� V�  CD1     SYS           ��:!� օ  FORMAT  COM           �2�� �Y  MOUSE   COM            0j� X�  �BR     ASM           ��V� B                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  �5                                                                                                                                                                                                                                                                            ��                                     .�#.�./.�-.�61.�33Ɏ����6x �z �"� ���x "�z �|.��|.�7�|.�+�|.��|.��|.��|.��|.�'�>&|)u.�%�|.��� u� |.�'�"|.�)�3�������3ێۋ� �� �RPu�Lu	�иJ�/�±.���B+�.�5����B+�����8PˌȎм3��ء|3ۊ|��.�.�..�).�'.+�� .���+Ã� �|���+Ã� 3Ɋ|P��3���.�X��=�r.�.�HH.�� .�67�� t\2�P.�#.�	.�%.�.�&7.	.� �HH3�.�7��.	.XP.�&� �3���.�7.�� X@@.H.�&-��ȸp �؎���3��.�>!2�.�7.�.�6�.�.�.�>0�t@3�- 2�.�7��.#.%.�	.�.�>!.�6�p ���% X.�&.!�.�./.�-.�#.�%�  p � Q.�	.�P��3�.�6+.�X.�6+.�++ڋ�.96s.�6��.�P��3�.�6.�X.�6����
��̋�.�-�ƴPW�_XYs��2�Q.�-W�_YIt�{��� 2�.)t.	.� 3ۊ�.�����R��.�5��.�0�.�.�>.uH�����R3��Z Zu&�.�FR3��I Z&�  .�.��&�.� u%�����=�s�R3����� ��� Z&�=��s.�0 �PVW��.���.;t4.�R3�...�� .�	.�.� 3���Z.�I;ы�_^X��^� 2��3ێ��1�x ��D��
�t������
Non-System disk or disk error
Replace and press any key when ready
 ��  �p                          5 p �� CON     G p  ��!AUX     Y p ���PRN     k p ��9CLOCK$  { p ��>�    � p  ��!COM1    � p ���LPT1    � p ���LPT2           � p ���LPT3    � p  ��'COM2    � p  ��-COM3    ��p  ��3COM4                        Np  �           	             P̀@ 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 �p    � @ h  	               (   � h� 	                �����NO NAME         FAT12    p   � @ h  	               (   � h� 	                �����NO NAME         FAT12    zp    � @ h  	               (   � h� 	                �����NO NAME         FAT12    ��p    � @ h  	               (   � h� 	                �����NO NAME         FAT12    	p�  P P P P     P�p .p  FAT12    FAT16    NO NAME                     $                   	  
                                               !  "  #  $                                                                                                               �����  ��������	����
��������������������p����r����s����t����v����w����T��                                                       ; Z x � � � � 0N   C ����K�.� �.� .� ��@ � �; �   �4 �  �- � �& � � 0 � 0� 0� 0� G� �.�>  tP.� .9 Xu.�.��c ��PVWUS�� �[]_^X�.�>  t�V u�E .� �.��.� � � �.�� .� �.�>  t�! u� �ː ���   � t�PS�.� [X�QVW.�6�.�>�� �_^Y�PS�.� [X�� � � ��������������>@ t"�A� ������ح���t=��t��������>  t�0 �=SOt.�.P�@ �ؠ $<u�>  t� X�.�.PQW�D������� � 3��_YX�.�.����             �p   P   P   p                  WSP3��ǻ ���/���t��PW� �X[_����s   NO NAME     NO NAME     ���  P     �                  (                                �   NO NAME         FAT12    ��  P     �                  (                                �   NO NAME         FAT12    ��  P     �                  (                                �   NO NAME         FAT12    ��  P     �                  (                                �   NO NAME         FAT12    ��  P     �                  (                                �   NO NAME         FAT12    ��  P     �                  (                                �   NO NAME         FAT12    ��  P     �                  (                                �   NO NAME         FAT12    ��  P     �                  (                                �   NO NAME         FAT12    ��  P     �                  (                                �   NO NAME         FAT12    ��  P     �                  (                                �   NO NAME         FAT12    ��  P     �                  (                                �   NO NAME         FAT12    ��  P     �                  (                                �   NO NAME         FAT12    ��  P     �                  (                                �   NO NAME         FAT12    ��  P     �                  (                                �   NO NAME         FAT12    ��  P     �                  (                                �   NO NAME         FAT12    ��  P     �                  (                                �   NO NAME         FAT12    ��  P     �                  (                                �   NO NAME         FAT12    ��  P     �                  (                                �   NO NAME         FAT12    ��  P     �                  (                                �   NO NAME         FAT12    ��  P     �                  (                                �   NO NAME         FAT12    ��  P     �                  (                                �   NO NAME         FAT12    ��  P     �                  (                                �   NO NAME         FAT12    ��  P     �                  (                                �   NO NAME         FAT12    ��  P     �                  (                                �   NO NAME         FAT12    ��  P     �                  (                                �   NO NAME         FAT12     ���r
��t
��
t.�.SQRWP�@ ���t  ��:u r�t � S����Î�[���� rXP� ����k X�&t 
�t�_ZY[� �C �H  ��t�H "��$?�D �.E �����F ������
���G S�\ &�G���B &�G[�&v ���
��&v Ë��@ u5�B u/� ����m����H t�1 r� ����l��) u�C u��he��/ �he��. �he��. �he���. �he���. �he��i/ ���w.�.���r�P�@ ��X�.��  .�6�.�>��s.��.��P�.��.�� .�.��3�.������.�����. �.��.�>�nv&.��.�.�n� .�>�mv.��.�.�m��.��3�3�.����� �Ê;�vF+���.����.�6�.��.���.���.���.���.���Q�
���
�Y������� ��6���� �����.�PQR2��ZYXPSQR.�� ��s� �.����6���.�� �Irw.�� �� rk.��  � ����>�ud -P ���ܘ����.���Ø�t�m��.���>�v.����2�I.���2�I����.�.�6�ZY[X�3�3��8��r�.����6��� � r�� r�� �.����6�����à�� ����� ����� ����� ��Ê�$����
À>� w5t�>�r,�>��r%�>��w�>�w�>� v�>�1w	�>� v���À>�$w�>�Yw	�>�Yw���ù �����%�<
w�����������
wCIu����Ð             �   ��	(   @    p        �   ��     �       @     @     @       @ @   @ @ �   � @   �	    01/10/84 �  p �� 	          �  � `	�           �  p �� 	          �  � ��	 $          �p���������� .�6�.�6�U� �P3���X.��.��QW�s�ؾ?W�
�t	�� ���� � .������������������_Y.�.�� .�.�� �L t�N �T J�V �d ��f ��� u6PSQRW�� �r.��_ZY[Xr.�>� t.�����.��� �
����% u@.�x @���u3�3���Ҽ �Q��P���r�� u&�G.�>&�G.�?������&� .�>� � .�>> u�f� t
��P�P�t��	��	��|	2��w	��j	��e	2��`	3Ҏڎ�3��4�����l ��n �� b�� � ����������������� ��,.�&.�>>�r�+�"�����Y.��PS3ێۋ� �� �RPu�Lu	�иJ�/��[-@ .��-@ .��X�s���u# �w�������s

�s��3��ء> &;�v= �u
�< ��> 3Ɏي���t.��.���	�  	X2�u �%��^� ��؁>��COu�>��MPu�>��AQu� ��r��@��������r�]2��,	��>�u�=�=����:u r�3ɋ=� ��(WRQ��rx�� u�'�	����ň6���?���.�:,v�,YZ_��r��u���w �>�(u�>�	vT��P�>�Pu��	�>�$t@�>�t�>�	u޶�.��*YZ_��r��u���w ��P��:,v�,�� ���>x u�π� 3����E6���E4�M#�u"�U�}���]%�>x u�x ��	M#�=������������6]
�t[��R�>`�u � �Sr��s��Z����u����6]���RS�>`�u �*r�s	�[Z����[Z����uـ>%v��>`��	u�	�>w  u����>>�u#�>] t�� ��ƾf����	 �u����K� ���&�>��COuK&�>��MPuB&�>��AQu9&�����=68w.r&�����=80w!r&�����=40s�-��>� �� +���>�u�>�� �.�>� ���W�A�&�=��_r�y 3��؉>����
��������������p �> �����������3�&�&��&�������].���]&���M�E&)��E&�2�3��ߋ:�s��&�s�.��@u�������r��I�is.�>�}�t	�=���u��P��E�=�����u�.�>�=.�&%���=�E����u�.��<r .*%r�.u .�����s�ߢ��.����� �2�� �r	&�>�U�t��WS�]�U�M#�E"�� ��R���ƈuZrc��?�MR��ZrV��&�G��t&�?t&�?t&�?u
�t:�΃���uػ�&�G��u&�?t&�?t&�?u
�t�΃���u����.��&�G&�W- �� &G&W
s���&�G�E&�G�E&�W
&�G�U�E�� w=@ r��U�E3ۊ]P��3���.�)X�����3ۊ]P3�.�)��.�)X��.�>) w|= ww�}GuEI���̀��
̊��.���N���NSP.�?�t.�?�u).��u"�Y.�G
$�<�u.�? u.�G
�t��s�tX[�6X[.�2.u.�
0u�/����"��.�0.u.�G,1$�t�.�3.r�u.�
1r�.�>t)uW.�>^ uOW�Y��.�| u#.�| u.�| u�E.�D�E.�D�E.�D� �_�Q���S�Y3�.�D�u.�D.�T���t�E�U�E�U.�\�]	+Ã� .�\�]��+Ã� .�\�]���+Ã� 3�.�L�MP��3���.�)X��.�>) w=�r��@�Q�,�� .���� �M# �U�E�.;rw.;Dv��
��L�.�L.�T�U�U�E�m��@u3ۊ�K���C�������ށ����}�=�R�U��+�Z�� - �� ��}Ã� - �� ��E���]�����U�E�� w�} wEr�E�E�E  ���]�[_�PRV.�>t)t1.�10u.�
0u"�Y.�| t.�D.Dsu.�L�m�] ^ZX�   3��>W&�]"��u>3�&�E�u&�U&�ERP&�E&�e��XZP��3���.�)X���t@&�E%�u�V.�>�tT��u@3ҋE%�e6�e4�E/H�=�r��������t�E-� �U).�&�!.�6�!3�.�6�!@�E2�����0�}'� �_&�=���t�L�Ø�д�Ø�а�� �Ê6]�� t1��R�\����3��ƣb��?���d�\�'�r�	 Z����u�Á��&�?t����u��|� sw�>`�EG �M#�E"�� �b�E�d�E�\�E�u �E&�
 w&�@r;��&�w�������&�W�UI&�O&�w�\� ��r���
 r�A �s��WS&�?t&�?t&�?t����u��[_����>u r�s��&���VS�6�<�t�4���<�\����]�]�6^��^�u �`d[^�PQRU3�3�3Ҵ��� u�� u��tE� @����.��� V����6��^]ZYX�P.�>>�u%.�>?t.�>?s���&�0 ��� $���" XÜ�SP��p��q��X$��p��q��[� �ϜP�P��p����qX$��p��qX����QW.����HH��.�.�PS.�6��ދ�.��@u>���R3��~ Z�u�.��FR3��l Z�  .��.��[S��s��������؁���R3���� �? Z�^X+���u.��SRP.��.��Z.�+����[_.�������Y�PQWV��.����WP.������X&E	_.;�t*.��R.�+  �й .��3����O�Z.��I;ы�^_YX�                                                              p .�0 ��� �GG���VPQRWUS��v.�0 �D�! �&��4� &�G&�g&�O&�W���u�+  ���u&�W�+&�W�&�G.:s,����&��.�Tr�.�0 � �G[]_ZYX^����	 ��       �� &)O���� ���� \��	������� ���Q������������������� 5�lttU
���� 5������� ����Ê&�2�� 
�u*��t�= ru���>� t<�u
�t2��
�u�& à 
�uM�&��u�>y  t� &�G t� A2������u�&����= ru���>� t<�u�� t� � &�G����&�G�)�����  ��t�2���������.� �7 u&�2��/ t���u	��  ���tKu���G�����
 u��Āu��j���! �P��0��0Xu��߀���(t
�	�� u��ð��Ë�QS2����㋏�[��u�Ā��Yt&�2���u����Y���> &�}t��&�E&�}2����㋏�<et<Eu�&����&����> &�}u&�E<et<Eu��������{ 2��
�u� ����ô�> ��u�X2�����U �
�u�" ��t� t�������s�� � t��� t��ô�! ��� � ���&�G�����Āt�
�N����Ë! �� ð<�� ��p����Ȱd��ȃ� � ˃� ������ђ����� �� ��ȵ �Ę�����&�P�>� t&&�E���&�E���&�E��� ����&�M&�U���������>� t
��������N �6���������������������3���ӹ� ���dr��d����в �ҹ< ������P�ƫX��ë��2���>� u2���
�t��� B��� W=XXIAXX� 
1XXXkXXX$B��>&8Et	&�=���u������� &�E$t&�e#����&�E#t����,&�E#u%3��>w  t
��r6�Uu� �&:Eu�( �N� &�w�y�>w  t��������þ � �&�EG+�&�EI�u�u��>r����$vN���&�%�?�&�E#u#�7 �
�\ r��>
�
 t
�>w  t������� &�g&�&�O��W3�&�MW&�MY� ���K�&�E@�u�� ���_�&�E#t� QRS� r	�u�� �\� �ar��>w  t��&�}"u���uz����  �� �� �� �)���r`��@�@���u���Ã�(��tɷp����&�u&�}&�M&�e&�E&�]&�U&�E  &�E  &�E  [ZY��
 �>���
 ���� � �� rK3ۀ>Nit�>N�t�>N�u1�>P�u*�c$�<�u!�c<�t�u�>V3.u�>X2s�[�C��Ê6[�>_�a�&c�d�f�h�>
u� r�
�>w u�'�À>t)u.Q�u&�MW�w&�MYWV� �y��K� �����^_Y���ö � � r�'�U� &�U�N��sL�tD&�E#u�>8 uP�6-�D	�D	�*X����>8 uP�*�6-�D	X�s뷲���v �&�mF���]À>w  t���&�E �À>w  t��&�}  t&�M ����&�E#u�ô��� ��  � s���� ��PS&�]#��!us��tn&�EW�>&8EuS� &�]#tK&0]#_&]#�>z u&�} u>&�E� &��.�>x uP&�E��� &�:�Xt���&�=���u��_[Xð����� �ߌ7���&�E���&�E$uމ"�&5��3�у� &�} t�� u�&;Uw��6+&;urw�&;Uw��+&E&U�-� &�6x �6-�/&�E#u����>w  t���J ��3�&�u�)�-&�u�1&�MP3ҡ)��)X��>) w= w�2�3�"� �M �� �&�E��>8 u:�,�6-�D�D
�d�&�&+�6-&�}"u��D
2����D	�'��(�&�E#u/����>8 u#P�6-�+&�D�'�&&&�D	&�D&�d
X���t�&�E#t�/�t�) 3��&�M��*12�;�s��PQ��� YX+�������� � &�E#t��t� �.2�.4�& P�3&�E#t&�}Gu&UI����
61�ʆ�62&�U&�}"t�>v �t
��t��t�V�� r��v &�mF�> tRX&�E#t�/�u0��?2�)"Ȉ1&:Mv�1�62��&:ur2��3�62��:v u&:mFt��u �XP�� s���u�4t��X�>�S�2��>w  t�f�>6u� �6 � t &�E#u���t���t
�4 X���� ���M ���"�&5�X��>8 uP�(�6-&�D	X� �6-&�D	�&�E�u�7��7�����Q�ĢD�	 �<򮊅 Y��P�t�&;UGu&;MIt� &�UG&�MI�X����tM�
�� �������i���������`@aAbBfFgGh�i�� &�&�Gu%�<� u�O$�,@.:w���F�.�.�0 ���Z�.�� �_&�E"�G&�E#% �G&�E%�G2��G�u'�t.�0 ���'�r�u�� ���� �_&�M#@�u|�G&�E"�G&�E%�G.�0 �>w  u%��% &�M#�����&�E#�G.�0 �7&�M#� W�u&�E# t&�e#�� �}'�&�M#� �}�w�.�0 ��_�O&.�0 �9&�e#��t&�M#��?w��;�w(.�0 GG���������ð��� �_�t.�0 �A���&�}"u.�0 � �O�W�.�0 t�� �<t<u�gR�Z�J��£9�8��;�9������ Q�;�9��7�YrQS3ۉ7�9���y[Ys)�Z�9PQR�<u�GZYX��9��u���u��9 �� �_�O�G�W�� �3�2�9��t#��
�u.��
�u(��&�E# t�/� t�63�3ۉ7�? �6 ô��� �� � &�_&�G�3&�G�2&�G&�O&�_	�7�&5�9��>8tPQ��YX�;����� &�E# t��QRFF��1&�E# t�/� t�"����ZY�ìPVP�&,�6-�D�dX�£"���^X� �ZYⳀ>8t�h��À�w��ðÊȸ� ��À>9t&�E#� tL&�e#��9 �;P�&�}"t&�}"t����>7 u��;TV� �6x �D	^�&�U�&�e�&7�QR�>9t&2��>8u� V� &�6x �6-�/&�D	^&�M%I�����͆�&
M&�UVW��r3�>9t%� &�6x �6:�<� &�>x &�z �82��9���t	���t�����_^ZY�P�>8u�92���v �X�SV�8u6P&�}"�� &�6x �6-�/�7&�D�;&�D&�D	�u&�D
X�9��&�U�68�7�^[���&�E�>&8Eu&�E#  u&�=�����z ���z  2�&�E# t&�M��� �O��P2��9�8
�tV�6:.�0 &� &�6x &�z ^X��� &�E� �} r&�>c�r�>t)u�> &��u��� ��ð���i &�E��� R�B Zr>�>c�r4�>t)u-W�u�6 �t��� �_�?���� �
 ��ð��WS�N3҉+� ��[_�&�U
�x"&�E# u�>w u�$t��sS�@ ��[�� �_� &�E# u���G�� �_&�e#��� u&�M# �� &�G<u� �`���u� � ����� �_�  &�U2�� �r���<t
<t<	u�G�À�2t���1t����� ��t��t;��ty��Ju� �P��.�0 �6� �6� �6�6�� �� ��[ZX�<�s�
�u����<t<t$.�0 � � �p .�0 ����.�0 �>�.�0 <t<u%�� u�&� ��� u���������<u�K ����Ë����tC�<u3������- ���t!��;�v�����>�������u�����x��u�.�0 �>����u�>� t���>���Q� �� �w
�� �w�Y����Y�PSW�p rb&�E# tZ&�]��%? ;�vM��
�u���Ȁ��
�2�@ƀ� &;Ev6R3�&�]���u���tH��Z�ϊ�����?����������
��_[XÊ������>&8Ut	&�=���u��Ê� 2�
�t�� �� ���p ��� Ð @ �>w  tYS�@�M[�O��xRPQ�ʰ���1YXtBS.��ڀ� &��[�.�> t�> u-P���p X�".�0 � ��t��>1 u���p ��>>�tŝr!� s���u
�x�>w  tS�@ ��[��߀�	t~��uۀ>8tԀ> u�2䚗p � 2�<t�SQR�  �����p s��	t��u� 3��  t	���������ZY[�S�N���p [s��u�VW���N�!�_^�ơ ���r;��t<��tHw/RQSPU�����������Ӂ��s� �*�:�r6�v	���� �	���S�N��p [��SVW��N��_^�݋VQW�5�&�M&�E# _��t�?*�Y:�sP�����P�%�r~X(f���:�t
*����ڊv	S�f��u%VW�NW���K�[_^��V�Z����r:�"S�N��V�C����[r"VW���N��_^[��A�F���t	�V������][[YZr�2��U� �&u ���w���4&�E8Du�&]#\#&�e#ߊ\#��&]#�<�u،D�<&���&�E4:,v�,���t��p QR&�U���+ɸ J�/At��A.����S.��).�
�u��<�2��[ZY�
Insert diskette for drive A: and press any key when ready

 &�}  ��?�3��Zt/�Hu+PR&�U��ZXr� �&8]tPQR��ZYX�t3����r��- s�����t�t��r� r�y� �v��^����x(�>t)t(�� t�3��>^ t�� r����uF�� ������P�u&;EWu�w&;EYu3�X��X�����ڀ�u��5�t��"�r��r	�xE�� ����� � ��þ � ��K�8��K�@�&�E# t1&�}"t*���u%&�}"t&�}"	t���`	����0������W�>&8Uu&	]#&�=���u�_�&�E#@ �&�e#��&�E# �RP���t� r
� ����XZ�ZZ�  RQSPW�	� 	� �_&�E&�M��&E	.��&�E����Q.��&�M3���B��3�&�u�����rD� ��? t7�?�t�Gu�� ��Y.����3��Y��W�	� �2��3�_X�[YZ�Y��^^��WVQ�	��K� ��Y^_�WQ�	��K� ��Y_�P3��&:EtNX�                    H H     P� ���&�>���u�b��tX.�. X�     �8     �� �� A     �� N �    KB �       �� Y ��    KB �       �� q ��    KB �       � � ��    KB �       � � ��    KB �       �{ � ��    KB �       �c � ��    KB �       �K � ��    KB �       �3 ��    KB �       � ��    KB �       � 1�PU.�
 .�. �&�F < uQ.�. &�f&�V��&�n&9F uD���ŋ�n�ЌĎ�.�n �.�^ ��&�n &�V&�f&�F  .�. ]X���<t&�F � �.;. r��&�F ��.�. &�~  u�&�F < t<t&�F .;. t������ ��؀>���u��r����!桌Ύ޾;P�p ����Xt��p �<$t�������

Internal stack overflow
System halted
$�                           2 � 	 �         ��           A:\          
$  �     �Qs�s�s                                                                                                                       �s�s�s                                                    �    �  �p                                                                                                                                 ���r�� u&�G.��&�G.���.� ��ؠ��.���� u2ɴ� �r�� t

�u.���3���.��I3ێ�&�� &�� &�RPu&�Lu��R�J�/X��;�t.��I�pY�+ȁ� 
�p�+Ȏ��pY�����P˸p �،����pY�z�����3���.�s� P�.�s� .�q�W.)s�� 
��.���ؾ0 ���p+�����.��.�>�.�6u.����Ȏм2�.�q.��.��.��.�}&�.�m&�E.�o&�E.�y&�E.�{.�s.�.�>� tR����H�!�H�!��.+���H�شJ�!����H�!�H�!H��&�  &� RP&�
 L &�   &�   �I�!.�>m����r&�EE�t�&�E .��.��&�EC�S3�3�P��X% �= �t� �P��X% �tCC��[�= u&�ED&�E .����- .����������A+�.��W��-� .��.��&�}&�E  &�  &�M��3���&�&�E&�E� &�E  &�E  _��.����p ���˃���3����� �&�6 �P�!�lP�$%�!�>� t�Y�sI.��
�t�ʴ�!+��ءl.��.���.����4�u9.�h.�d.+h�J�!��H��&�  &� SD��& @.�6m&�D��	�I.�h�!�.�>l t.�s3�.�}�3��� .�s.�}�0�  .��.����3�3.������6�j�R7�p ��&�� .�� t.����.�>l�u�I.�>l t�j.�U.�h�I�!.�� t%S.�^.�`�J�!��H��&�  &� SD[.�>l t���� �Cs��R�D��D��Q� A��Q���PQR����H�!�H�!rk���I�!����ȋ����+؃�+�rK� =��!rs�؀>MQ u�5� �?�!�>5�uY�>8fuR3�3ҸB��!rF �� ����� ;�r��V�G�<�>�!��Z�������O�O�O� K��!R�>�Q t�>MQ t�V�GZ��!A�о�Q�>MQ u� ��< uT��Q�< uL��Q�< uDR��X�GZ��!R�>�!�OQ� ƇPQ�NQ�
�!��U��FZ�OQ
�t��MQƇPQ ��Q �5�MQ �PQ��D� �
�u���Q�|:u�T��
�u��E���R �C�ZC������H�!�H�!.�h.�d�HMA not available: Loading DOS low
$Fatal Error: Cannot allocate Memory for DOS
$�% r��	��	�!� �F .�s3�.�}.�l �� r.�s3�.�}.�l���� r������ .���9 ����M ���	 .���$ �.���0 ���p+����W��.��.��_�W.�6q�[.�q+��[+�.�søp-0 .� �ۋ�t�H�!rQ- ��&�!  &�( SC�WQR.�>mOO�&� ;�r'&�  ��É�؈  �   +ˉ ��- ZY_���	�	�!��p ���M uH�C�/� � ����� Ht	���=@ r&�� Hu�t�����&� 4&�> 4u���ø C�/<��PSQRVW.�>l�u��_^ZY[X�     �           VDISK  V3.3                 �       VDISK3.3�  @  �     @3��ءd .���f .���H� �!H��&�  &� SC@����d / �f �4 ��3����W������ �  ���_�                ��   �  ��  �                                                  �d�u.�>��t	.�>��	u��ȋб������� .�h.�j� �V���Ìø��+Ã������+��p �؉>�� ��3��؎N � � ���t����ؾ ��� �������3Ɏپ� �� � �������������>m&�M 2�&�M!���X����6�+�&�u��&�E  &�5��3�.����\ .���.��3�Q�? ���t.�>�u�<w��Y���Y�Y�| t� @��ƫ�ث������� �� �����.��A�.�6m�4,A:t�t���u���p �؃>/ u�/� .��.���U?.��,vRP�F�=	X2�.�b.�d.�>m�}��U.�>b&���&�E�;���.b� .b.���?�3����>�X��.��2�.�b.�d.�>m�]�U.��2��]�>b&���&�E�;����b� b���>��AQ�; ��&�E�  &�E�  &�E�  Y��>��t� ��  �� P.�.m&�n &�^ �øD�!�u63�&�^ �ú�S�D�`�!r!��S��S3ҹ �����u=�v�� �&�~�t&�n뮁>�  v"�� �>� @v��
 �>� �v�� X.�m.���G?.���GA�_��=�B�S�[[.�>� t-�=.�b�O.�d�O.���O
� ��.�b.���=�=P�L �uX.�>m&�M .:�s.��2�&�M!.�d&�E.�b&�E���X���X.d.���<=&�5&�}�B��>��t�>� u�>��sq���tj�=�S��d��3�3��i�b��<��p ���� ��.�b.����.�d.����� .�.�&�����.d.���<����2��3۴>�!� �>�!C����P��=��!s� ?�P� �>�!X�شE�!�E�!��P��6?��P��.?PSR�����B�B�B�B�B� ���&�>���t���r&�G@t�����B�B�BB�B�Z[XP�d+h�`�T�X�>d�ǉ>�3��>����� b.����;���w������;�d�h�^��+شJ�!��H��&�  &� SD����H�!�H�!�d�b  ����+�KK�J�!����H�!�H�!�h�d�I�!�V��3��.�� ���< t���&�<
t��G��.���� u.��.�    �ȋ�.�>� t.��.�B.�F.�J.�N�` &��3��K�B.�.�^sV�=^� ���������.�b .�&d �!.�b .�&d r� &9�t�	�f �!���&�.�&����3�3�&����tFF���2�pY+���&FF���    
Memory allocation error $2��V t��?�G�G  ��.��W�e ����.+>�Y&���&�M
�t�G.�d�G  �G.��- .b.���:�SR.��.�&� %���ظJ�/���u�  .�dZ[�.�6�&�E.��.�&�&�E� &�E  &�E  �PSQRWVU.��&� ��&� .��&� .��&�
 &�. &�. � &� ���&� �؃�&�> &� ���3��
 �� &�F  &�F&�F&�F &�^&�/���߃��. �. � ��؀>���u��r3����� �B� � ���  �G�8 �< ���$ �L�A �E ����j�N �R ��( &�Z�� t1�?�t,�KBt�� �uR� ���&;�Zt�Q�Y �W �j��, &�Z�� t1�?�t,�KBt�� �uR� ���&;�Zt�V�q �o �*��0 &�Z�� t1�?�t,�KBt�� �uR� ���&;�Zt�[�� �� ����4 &�Z�� t1�?�t,�KBt�� �uR� ���&;�Zt�`�� �� ���8 &�Z�� t1�?�t,�KBt�� �uR� ���&;�Zt�e�� �� �j���&�Z�� t1�?�t,�KBt�� �uR� ���&;�Zt�o�� �� �*���&�Z�� t1�?�t,�KBt�� �uR� ���&;�Zt�t�� �� �� ���&�Z�� t1�?�t,�KBt�� �uR� ���&;�Zt�y��� � ���&�Z�� t1�?�t,�KBt�� �uR� ���&;�Zt�~���j ���&�Z�� t1�?�t,�KBt�� �uR� ���&;�Zt���1�/�* �� ��؀>���u�'�r��p ���@]^_ZY[X�&��&�D�G�p ��&��&�D�E&�&�\�Q.�d.����&�  A&� Y.�d�                                                                                                                                                                       �    []|<>+=;" .��  �.��.��  .��  .��  .�8[].�:|<.�<>+.�>=;��s���S&�&:s� [�#.�6�SWU��.�� uC��_r<��t7��u.�� u��&.��AtN�.�<=u.��C�HsŬ.�C�N.�6�.� .��&��6�.�</t6.�<"t.��uT&�G2�.9�s.����CC�&�� �i.�� �`&�G2�@���&�2��tCS&��� [sACC��.�� �4&�G2�@���&�2���@�&�2��tCS&��] [sCC��.�� ]_[.��.��.�6�.��.����P&�� u.��.�< u� u	.�� �P���� X��X���UQ&�O2��t�o	��s� ����.�.��Y]�&�~  tE��E�.�����rJ.�&��P.��+�.�X.�6�.�< u&.�|�:u	.��	 �&�? t&� u.�� �	� ����
P���� X��W&�.�>�&�&�eP.��&�EX<u
&�U&�M�Z<u&�U�P<t�<t�<u&�U�><u.��@&�E&�]�+&�u&�MP&�Gt��	&�Gt��� X&�Gt� _�.�A P&��uPSRW.��	 ����[�_Z[X���o�� �t.��  �&.�>�	uW� @t.��  �� .�>�	u@� t.��  ��.�>�	u&� t.��  ��.�>�	u�  t
.��  ��.�>Au.�>� u.��	 X�PV.�
�t<:u.�| u.� �	�TsFF��^X�VR��.��Ar
�t� .��FF��Z^�<�s<ar<<zw8$��4SW�>3.8tPQR�e�»��� ����!ZYX.�].�ECC,�&�_[�P.���.�&��.�<+t
<-u.��F� X�PQRV3�3�S.�
�tB�� r92�������� r,�ڋ������� r����� r��� rՃ� � rF�[� [.��t
���҃��� &�w&�< u����t�F&�< t`F.���u&;Lr6w&;Tr.&;Lw(r:&;Tw �2&;L|&;T|&;L
|&;T���	��u�.�� �����&�$�.��	 ����.�^ZYXÜ.��u�Ýp����<0r<9w,0����PSRW&�&�
�u���L<u?G&��	��@�&����@�&�GG&�-�2 s����u�.�� ���&�e��&��.��	 �����_Z[X�PURV�.��<r<��.��t<=u&�~ uq�.��t<:u
&�~  u\F�\&:F u
�tRFE�&:F uEF.�E&:F u:FE�.��@t&�G  t&�~  t"&� t<:u	&�~  u�< u&�~ :t��.�6��^Z]X�PWV.�>�.�
�t�_ u$.�A^.� _�?^.� _&� u2.�� �)XV.�
�t�- t�\sGFGF��.��.� G.�>�^_X� t	P�����X�SQ�8�	 .:tC��AY[�PR.�
�t8�r,.�|:t&� t.�| u <ar<zw,`�д���?��.��	 ZXì�" t�S u.�� t�.��At	N����N���SQ<t-< t)<
t%&�}r3�&�]��&�9 t3�&�	C&:t��<Y[�SQ.�� .�&��< t6<	t2<,t1< u�< u� F:��&�}r3�&�M�t� C&:t��< Y[�.��.��u.�� :���.�;�t
</u����</u.��@��VS.�>� u'PQRWU3��޸ c�!���]_ZYXt).�6�.��.�6�.���< t:r:Dw��FF���[^È ;� � �   �  � �     c   �  � �             � � /X               � ;�       � �    � � ON OFF  � ;	!!&!   �  � !    �  �  � !   � �      8!;>!   �  � G!    �    X!;`!t!   �  � i!    �    �  � }!     �     �!;�!   � �   �!;�!�!   �  � �!     @    �  � �!            �!;�!      � �   �!;   """$"0"     � � /K     � � /N     � � /F     � � /T     � � /W    D";L"L"      � ^"     � ^"   n"s"w"{"HIGH LOW UMB NOUMB                                                                                              PROTMAN$         � 7�!��Q��Q��P� =��!s	� ��Ë�3�3ҸB�!�V3Ҹ B�!���V���P�+�J��+Ѓ������ڎ�3�.�V�?��!�PWQ�����uO���
�+�.�>VY_XP�>�!X�r;�t,��P�,��>�
s��6��6X�6V3��6Z�6��3
��~�+
r����� �� <
tL��$�>� t(P�
���
�ģ�X�>�r�� t�>�r&�����	s�>�s��	�')���	��>� u��>�t�>�t��Ht
��Iu���ɀ�Wum��뽀�Iu
�U'rB��뮀�Wu8�F'r3� X�!��S�ˀ �X�!�X�!2�P�X� �!�q�X[�![�X�!�q���Yt
��Zt��0u�Z�V�W���Buc��&r^��  �� 3ɋ��s���E=��t�>� � u��� ��u�� ��� �Ճ>� cv���   ��� ���� �����������Cu=�&r8�� 3ɋ��Bs�|�$=��t�>� u�� ���  �ܴ3��� �!����Mu{�E&rv��!3ɋ�� s�:�7=��t�>� u��!���! ���p ��.�>�! u�/ ��/� �X���Ht�����%r��?"3ɋ��s���
=��t�e���-���Uu|��%rw���}s.�6�.�����.��"�u�	s.�6�.������V&�<t<
t��&tF��.��"&� ^��s.��" �6.��" .�>�" t(.��"� ��Dt�	�A%r�.��" .��"  .��" �6|�~�6�"��"�� ��&��rB��"��"��" t�<�t��"��t;�"}��"���v��"�"r9�"s��&��&�< s��#)�����r�V��VV.�6�"�D �u.�6m�| r
^^�� ^�9�.�>� u.�x  .��".�z.�m.��.�����G P� �V&� �P&X.�m�G �%.�x.��".�z.��"�=.�>�" t�.�>l�u��^� �$��V�(�d^.�>� t
�<.��  �:�.��".;�"v^���.��"��.�>m�D� �t(.���r�� t&�U&�]� t&�U&�]
� .�w
�t��D
. ���Ȋ�&�U �����v�k�.����r�& E . �.�|.�.m&�n &�~�t&�n��.��"&�F.��"&�F.�.�".��"!�c&�F��&�F��7CC&�V �S�!&�F.�>m&;Ev� R.��"&�V&�^ZB����{�.�>m&�M"&�U$.�6�"&�u"&�]$�.��"��T^@t.���2���.�� �&�A� ���.�>�" u=�J�  �/�u1�� �u.��"�. .��V.�d.��+ѻ .���U.��^�^��U��U�&����Qt�(�0"r�.� Q .�1!  �� 3ɋ���s�� .�/!���9=��t4.�>� u.�� ��u.�/!�.�1!�VW.�6� � Q�1&_^�.�>/!�u
�%���+V� .�> Q t� Q��Q� =��!rI.�\��.�/!.�1!.�d���.;�wH� Q�< uFF.�>yW����%_.�d��3��$s&���t�.�> Q t� Q��Q�%.������nV.����s�%�.�\�>�!��= u�+V��QV�%�dÀ�Fu0�!r+�3!3ɋ��s���=��t
.�� .�R!��.�R!.���6���Lu0�� r+��!3ɋ��s���=��t
.�� .��!��.��!.������Pu� r�r	�#�j������Kt� �{ r���!3ɋ��6s��V��$�� =��t.�� ��u.��!�.��!��.�>�! t.�>�!r.�>�! s.��!���.�>�! t.��!��.�>�!�u .��	 .��� .��  ��V�$�I�.��!.��.��!.��.�����5���Su^��rY.�MQ.��Q  �QQ�E���
�t< r,�G���Qr��!� ��Q��< r	�G��\Rr��ρ��Q.��Q� <
t�s��y���XuA�jr<�S!3ɋ��%s�_�(=��t.�� ��u.��!�.��!��.��!.��.�� ����1t� �!r���!3ɋ��� s��n=��t3.�>� 	"u.�<"��.�>� -"u.�="��.�>� 9"u�.�>"�.�><"�p ��u
�� ��.�="��.�>>" tS�R�!&�� [�����Vu�r
�s��� ���Nu�r��r��؀�Yu�Z�V�����0t����t��Z�V�N.�hH��& @.;�w.���.��.�6��  ��=  t=��u������U�"�_ ú�U�"�U �Z�RV��U�"�6����t��!F����U�f"�* ^Z�Q�V��6Z&��V�Z�Y������V�="� �� W�1"� �W���
 .��=
 r3����0�O��0����"_�2�.�� HtHtHt.��" �.��"��.�l �.�l��.���M t.�>�" t.��"� ��@ �ۋ .��"��� .��"��.�>�" .��" t�@ ��.��"� �V.�6�"��
��"� �^��b�!��.��� �PQW3�&��"&��"&��"&��"�&��"�� ��"� ��"�_YX�PSQR�O �\rA��3ҋ�B&�  &� �u&� ��&�  & ��&� ��&� ��& C��<Zu�� ZY[XøX�!&��"�X� �!�3���"�X�!�W��� t�</tN��+�$�<Su� &��"��<Lu�o � s�N�� NN�_ì<:uJ�rK���� rA�F �<;t��] t:�M t4</t0<,u!�� r�c� �! �<;t��8 t�( t</t� N�ø ��N��P��"��&��"X�< t<t<
�< t<=t<	�PSW2��&Ƈ�" &8�"u&��" _[X�<r��SWV�>�"�u��"
�t��2�� &���"
�t�^_[�SW�ٷ ��&���"_[�  .�>�0u��ar	��fw ��WÀ�Ar	��Fw��7À�0r	��9w��0���SQ�3�3�3�3�.��0
 &���r1
�u&�L��xt��Xu	.��0 FF&�F��r� r��r����N�Y[�P��.�&�0r��X��.�&�0���3��X�Q��蒱���Y�V�R�!&�� =��t���^�P&� = t=	 t�&� =SCX�QR�����r/��3Ɍ�;�s(���uA&�  <Zt��& @������& ;�s3�I��ZY�.�>�0u	��=��u@�PS�e�[X���"<�u���
�t���PQ��r7������&��"�) <�t 3�A��s���� r����� 
�u��YX���"�SV��"2仗"��Ë�^[�SV2仗"��Ë�^[�&��"�R��"���t���Z�P�z r!���t�( u�* &�  <Zt��& @����X�P��"
�X�&�  �&�  &� HI&�
 DD&� EN&�   �P&�   �  &� &�
 &� &� X�PQR2���;���3�;�t�H�uA&�  <Zt��& @�����ZYX�SQ���r93�3���t'�t�u&; ��&� &�  <Zt��& @���ԎË��u�Y[�P2������"
�X�SQ�،�&� �� ;�wE&�  &� &� &�  M�@����+�H&�  &�   &� �  &� &�
 &� &� ���Y[�SR����t+���@�r$P���W�[�t;�v�������t	�t�r���	���X�u3Ҋ��\��t����Z[�P��r��� u��&�  <Zt��& @����X�P&� = u"&� =FRu&�
 =OZu&� =ENu&� =  X�&�  &� FR&�
 OZ&� EN&�   �PQR�}�2������3���uA;�t���u��&�  <Zt��& @����ZYX�PS�E��
 ��T��[X�PS�R�!&�G���&�  <Zt��& C�����=��[X�2���"�X�!�P��"
�uX��� �  &��" � X��2���"�X�!�P�k r��� u�D &�  <Zt��& @����X�P&�> u"&� =HIu&�
 =DDu&� =ENu&� =  X�&�   �  &� &�
 &� &� �V�R�!&�� =��t���^øX�!
�u�X� �!�.�>�" t:.�>�"t������� ����r��A s��s r.��".��".�"�.��" .�d.��� .��".��".��"  .��"�.��".�".+�"�u��H.;�"����  � SD@.��".��".��"û��� H�!�tK.9�"wC� H�!rH�����3�.��".��".��"��WV��&�  D@&� P.�6|����<:u����<\u����
�u��� � �
�t<.t����� �X^_��ָ =�!r8�ظB3ɋ��!r$ �� ����t	.��"���������.��"��� >�!��.��".��".��"�ˎû�"��K�!Ü.��"��r.��" ��&�
�tF��.��"&��.��"��.�".��"  .��".9�"v��P.��".�>� u.;�"u.�>�" t��X��X��.��".��"H��@+��أ .�>�" t.��"�.�d.�b  �S��.��"  .�6�".��"�1 &�<SIu"&�|ZEu&�D�u��� r.��"�
 �ދ�[��[��&��buF���3�3�&���t9��
t4P���EXt�* r&� ������
�F�� �� ����u� ����������À�0r��9w��0À�Ar	��Fw��7���� r�? r�[ �����D�u-�R�!.��"�C�/.��".��".�>�" u�<r.��"�����P����.��"�t�.��"= u�X����.��"�� �؎�;�w&�>  Zt\���� ���A+����  M�  � � SC��&�  M&�   ��&� �C��C+�&�  M&�  &� &� SC�G& &�. &�  M��@+��؎�&�  M&�  &� &� SC��&�  Z&�   J&� �3�.��"&�� ����&9> t�" r��� r&9> u�&� A &����À>  Zt�� @���������rq������+��؃���&�  M&�  &� &� SC��&�  Z&�   J&� .��"�� &��$ &�3�&�=Zt��& @����&�. &�  M����.�>�" t$S.��".+�".��"� J�!��H��&�  [�.�>�" t!.��"&�$ &�>� �+�r;�t�����  Z�C:\DBLSPACE.BIN C:\DRVSPACE.BIN C:\DRVSPACE.INI     
 S.��" .��"  ��;� =�!r_�ش>�!��;� =�!r�ش>�!��;�G��;� =�!r�ش>�!��;�2�v;� =�!r�ش>�!�v;��t;� =�!r�ش>�!�t;���;��t;.�6�;.�6|.�~.�6�".��"�4�'��@ r.��"���.��".�"r.9�"s�B ��.��"�?��A r�.�x  .��".�z.��"&�,.�F ur.�� .��.��.����&�?�u'&_��&�?.u&�;u&�w&�.;�;w.��;�j.��;.��s�HY�	�!��t.���.���G �h.�x ��������.z.��".��"  � .��.��+�.;�"r.)�.��� .��.��".��".;�"�B w\.�6�".�>m��B �� .�w
�t?�D
2�Ȋ�&�U �����w$��r�& E .�|.�.m&�n &�~�t&�n��D ��C � .��"&�F.��"&�F.�.�".��"!��&�F��&�F��7CC&�V �S�!&�F.�>m&;E�E wU.��"&�F&�^������.�.�>m&�M"&�U$.�6�"&�u"&�]$��T���.��".��+Ѹ U� .��3��[øJ�  �/�uw�� �tq����J�/ .��".��" .��"  .��"P.��;.�|X.�~����.��".�".��".��"  .��"�2?3�� �� ���J����/�3��U�øJ�  �/�u:��,A��.�6m&�t�X�����2�VQR�J� �/ZY^:�u&�dC����X��������� �    DBLSBIN$ PSQR3ۊ U�ú�S�D���@�!�p ��.�U t.� U���1.��S:,v�,ZY[X���SP ��S��S  �U  �<t!<
t=< v</t��0�9 �Ur��r����U u���U% ��S��S  �� ��V�Z�����rQ$�<ArK<ZwG��U� ��U�u6� ���U؋ȩ� t ��r<:u��S.�� �.�� [� ��3��ÅUu3�� t� U�(��� t��S��t�� t��S���  t��T���T��3ۊ�S�� u��S( �㋷�U��S� ���U  t��T��S�U@ t��T��S��S���>�S�>�Sw=u$�߃>�Su	�>�SPu�$�>�S(u"�>�Su����>�S u���>�Su����S��S��S�&�S�&�S��S��.�V�'3���3�.�P �t��<
t< v���.�P ����QVW��M��R� ���F�E&�=;t0&�G$�F:D�����u�&�=t!&�=
t<[tP&�<?u	X��
�0��oXu�_^Y�_^Y�Z��y<
u�돪$.�T<[t[<Ot<Et<At<Jt�c�R<
t<t</t�(u��NA.�>TYtb.�>TDt4.�>TIt,.�>TWt$.�>TSt.�>T1t� �$tv���
t�� �th�� ��
t��tZ�� </t[���
t]< w��W�� < t�<	t�<=t�<t*<
t&.�R.�Q� < t<	t<t<
t.�S.�Q� <
u���&� G��&� G��&�E� <
t��� t��i �S
t���| t��Z �<"t>< w�.�>TUu<
t<u�&�E� �.�D?��<
t��.�>D?t&�E� �.�D? �!�.�>P t.�P �.�P��&�I�Y.�>V.�>X3�.�6Z���� ��.�>P u0.�>Qr(&�.8Ru.�>Qu&�D.8Su�&�FI<
u����Ru!+��ش�u���u�l.+�=% r�+۴��tCC��R��t>
�u:��bt��?u�wW�[��R���et��Bu#��W�D���R� ���R��t��r�����P+���&�.;<Wu�&��.;:W�u� X�QV+��XrL<[uC�@<Nu�u8��&�D�0�.<1u*�6<
t#</u��+$�:"u��R��:""u���R�����^Y��Ru���s��+ۿ�R�s@��R �QR� �������
��Pu���������
�:�u����RZY� ��R��R  ��R��&�R��g+��r.$<[t(<OtM<EtI<At<Rt�<Nt<0tn��ti��@�c����^�b�6�R�>�R u��rL�rG���$��Zr�Z��R�5��	s0���Bt�� �#B�ڈ��Rۉ��R���R���r��r�߉��R���i�
�u+��� +ۈ�R�>�R�tCSۋ��R�� �*[t	C:�Rv���R�>�R u
��Ru�� ��� ��@ ��&�N ��R&�b ��R��R�� �>�R+�&�J ��&�6� 
�u�6�R��6�R��W�
��Ru�>�R�6�R� ���>X��	������R� ��C:�Rv�� ����>�R���+X��	�9��U�	�6�R��R�w��R���u�+��� ���u	�V+�������ROuۋ��R�������'�ۋ��R��R�V+���+�S�=[r<PQVW��R��_^YXt�tW����_ru�^���Y�r$<[t�����Q� ��RG.��G���y .�6�R�u��R&���t�FG���
+�.�>�+�YQ�Y����F&�   �& �>�R t�@ ����R&�N ��R&�b �V�X�QV��+ɬ
��tn<�ti<
�tdA<=u� �$+�I+�&8t%��QV�^Yu'&�==u!����V����.��+��&�^��t��
t�	Q����Y���<t<
t���*��&�.�>�^Y��{ro$<[ti<J��u:&�D�0W��R�� t%��R�� t���e ��_uQ��VJ������^Y*��+_���$�G< r.�>� t	� �GG��r�G<
u�����P+�Q��V.�V+���rC;�r�^YX�PQ.�VV+��	 ����^YX���r"$<[t<Ju.���.��� v����W�r��%tG%��:�t��_Æ�������PQV���^YX�PSQRV��>�R�R��������0�&�R:�Ru��p����:�u��� ۋ��R�܊>�R�	� ��´��.	��´�� 	��´�&�G<	u� < r<$t�	���Ns����Z��^ZY[XÊ�R���7�D�>�R�tR�,�!����R*�Rs��R��R �� S�؊>�R��R������X�<�Ø�
���0����0��Z��[����!u�>�R�t�,�!��*���s�
�t� 6�R�P�����R<�tS� 
��R�P �[X
�uZ�!t�<Hu��v���R�����<Pu:�Rs��R��C�����c ���Ru�<Bu�6�R�^ �p�<?u��R���� �&<t<u����,0v�:�Rw¢�R�G���벷 ��0P< s� �д�!��U�FX�S0�
��R� �[�S��R��R���R��Rt� �� 
�P �����X�>�Ru��X��Z��[��S r�u�<t<
t�����< �\�r��t���<
t	�) r<
u��+�� r<0r<9wP�
 R��Z��X,0����Ã�r&���ù  ���Rt� ��Ru�P����Ru��u� V��X$tQ��+ۿ�R�
�t%G:t�y���M�� ��G���!���=��Vu� �!&�
�u� < ru&�< r�д�!�于X�� �
�u��?u�X��R�!$�:�Xt:�Xt�>� t�<uЀ�R��X�~�^:�XtX��X�0��PSQR������}�s�UW���!
�u��!��U�ZY[X���RtC��Ru<��R��R�D ��Q
�t'��Q� �ˀ���~w��Q���QA�g��'K���G��W�À>�Ru���Ru��R�Y �<t'<
t#<[t<]t</t< t< t<	t<=t<,t<;����r<
u����QV�ج<ar	<zw, �D���Vu<=t
<t<
t��^Y�P.�b��.d.�b  .�d.;�s#.��tV.�6���+�H&� .�&��^X�ú�V����.��".�"�.�6�".��"�j.��".��"�,0r<	w����S3����rJ�S�
 ��[À� r;����r/< t!<,t<	t.:�t</��t<
t<t
�u�.�V.�Z���[�.�� 3�[��WPR3�3Ҹ �PrMV�CQ� �^u=���<u5F��L� �*r'����wFFZX_;Du
�� t;Tt4FF������^Y_���T.�KQ�T
�L� �� r�FFWQV�D� r}�T�L� B��!rȺ � �?��!r�;�u��T�L� B��!r�V��^� ��
�?��!r�;�u��D��AA���w��6 <u&�u&�uWP.�KQ�DX�<u	_&�E&�E^Y_4FFI�� t�h��<u&�= tWPQ&���2��YX_�Q��J&�GG&8t&�=t�����)����<uG�&�}Y�P� B��!Yr	3�3��?��!�V�. r�FF���!A.� Q�Q�<\t</t�O� � Q^�P�<Ar�<Zw�|:u��Xä�|� u����V��U� &�
�t��!F���� .�>Ut���ô	�!�� s��P� Ë�3��D�!�u�>�!��=��!ð�MS DOS Version 6 (C)Copyright 1981-1994 Microsoft Corp Licensed Material - Property of Microsoft All rights reserved NUL CON AUX PRN \CONFIG.SYS A:\COUNTRY.SYS                                                     �COUNTRY   @\COMMAND.COM                                                    \COMMAND.COM /P \MSDOS\COMMAND.COM A:\MSDOS /P \DOS\COMMAND.COM 	A:\DOS /P  /P                                                                                                                                                                                                        �                                                   CONFIG= MENU COMMON [[BREAKCBUFFERSBCOMMENTYCOUNTRYQDEVICED
DEVICEHIGHUDOSHDRIVPARMPFCBSXFILESFINCLUDEJINSTALLIINSTALLHIGHW	LASTDRIVELSUBMENUO	MENUCOLORRMENUDEFAULTAMENUITEME
MULTITRACKMNUMLOCKNREM0SETVSHELLSSTACKSKSWITCHES1    P                                                                                                                                                                                                                                                                                                	      p �� 	            � `	�             p �� 	            � @�	             � ��	 $          UU5U5U5U5U5UNU5UgUFHSTDICN 
Unrecognized command in CONFIG.SYS
$
Bad command or parameters - $
Sector size too large in file $
Bad or missing $Command Interpreter 
Invalid country code or code page
$
Error in COUNTRY command
$
Insufficient memory for COUNTRY.SYS file
$
Configuration too large for memory
$
Too many block devices
$
Invalid STACK parameters
$
Incorrect order in CONFIG.SYS line $Error in CONFIG.SYS line $ONOFFStarting MS-DOS...

 Press any key to continue . . .
$MS-DOS is bypassing your CONFIG.SYS and AUTOEXEC.BAT files.
$MS-DOS will prompt you to confirm each CONFIG.SYS command.
$
 MS-DOS 6.22 Startup Menu
 ������������������������
$  Enter a choice: $F5=Bypass startup files F8=Confirm each line of CONFIG.SYS and AUTOEXEC.BAT [ ]$ [Y,N]?$YES$NO $Time remaining: $Enter correct name of Command Interpreter (eg, C:\COMMAND.COM)
$Process AUTOEXEC.BAT [Y,N]?$WARNING! Logical drives past Z: exist and will be ignored
$Wrong DBLSPACE.BIN version
$                                                                                                                                                                                                     �t|�=p   89:;<=>?@ABCDEFGHI	J	K
NOVWXZ[P\$!efhgl
Pi����T�T�U�U�UTKT�QR R�U�U�MxL�\�V�]s^%V�]�]�]�VDsLhL-M/MDDqMD�]�]9VV�L�N�]�]"M9HVHvH�HFJTLJ��sMR@YM�L+L�LMJ�`)`e`��+�:���9�����Ba[�{��_����_�ӡU��^>_�@�@eM�MAJ�N_��I��L�Ұٲ2�J�����D�@
M�@�J�Kx�^��O^�D���D|?0G.n�LGg��TC��/o����jkSk�H0P�0P�OP�(�w�����B��ήxIJlI�O��m���4DH�0PP�P+��P:��PQQ4Q9QDMS DOS Version 6 (C)Copyright 1981-1994 Microsoft Corp Licensed Material - Property of Microsoft All rights reserved <v���.��=PV�72��u��5Hu����+Hu����!= u�i �= u�� 2��> t��^X��.��=�0�.��=�0�.��=��
�2��.2��.��=��XX����P�6��6���$w܊�����lwҀ�3rt���dwt���Qt���bt���Pt�UWVRQSP��.��=������������3��r�0u�>�!�&����0�<��XP�&. �0 .��=����ӎۓ3�6��6�& 6�W6�L6�J@6�X������
�t��YtD��w6�>  u7��
�26�:6�#6�  6�"�P���*X6�X � 	6�7�tP�NX.���>6��6��6��6�&� ��.��=�>�  u'�!���&���F ��������X[YZ^_]ϋc ;0u��� �-S�.��=&��X[YZ^_]&�&�.��=&��UWVRQSP&�6�U��F]�.��=�6�� �@6�!���r&�F��s�6�  �Vr��nXVP����A�D: � ��*X^s�6�$2 ��P��.��=�
X��&.��=� 	�
�X���r=�&6����=�y3u��6�6��5�t2� ��B�u&�e6�������6��6�!&�&�&���P��.��=�
X��&.��=� 	�
�����r��6������c8�3�Pr�gs2�= t
��$��Xs��.�&�FC �t�$2 ��&�nE�.�������d��2��l � �}��L���2��2�6�$� ���V��6�>J t6�$S � ^�PS.��=�$�<�t	:�t������t�&&<�t�'�<�t�#[X�VQS�$��=���;.�<�t:�t��2��������2�.�:�t��2�[Y^ø .��=�#�����������u

�t���� ��t��t��u���t��Fu�� p .��=<u�7<u�� <u�<t��� t�w��  ��  ��
r� PSQRVW�� ���t"���؎���3���� ��� ��� t_^ZY[X�T�i @�1�l� �� � � �1����!_^ZYsRV��G�c ������!��^Z[XA�� �ش>�!���G1�_[X�0�R�ӻ��W�GZ� �� t� �>�u'�� PQVW�� ��3���� ��� �_^YX�&0 �& �o��uj�uA�"�\X���HR��It6ItLIt4It<IuC��H��&�=Du@&9Eu&�E� ��ȋ��3�3������� t�X �3���|������U��60N��&6 �VWQ.��=<u�����3�� � �Q�Y����<u�����3�� � �Q�Y���Y_^���.�6x?.�6z?PU��F]�E	��.��=ð�Ã��t*PR&�F&�V���t��2����ZXt%.��=���ËW.��=���O�_��PVR.��=�:�t��&�V �bZ^X�
Divide overflow
 You must have the file WINA20.386 in the root of your boot drive
to run Windows in Enhanced Mode
YNyn @M;S<>==?KRRAA[R}STTS�S�R�S�S�S�S�S�ST�	�W��G�_���.��H� �R�P�:��\��D6�Vð���r���ww
�t�
�t��w���} ���T�L2�ð���s���<s��<s��ds�QR��� 3ҋ�S�=�6. �6=[��=�����6. �"=2��.��=Q�  ������������
΋ѡQ�����Y
P���  VS��� 3ҋ��\=�6. ��<[^������;Tt�=6�s=�TVQR3ҹ����������Ⱦ�# ��s��� �$ ��� �QB�P� ZY^ô �;�r�+�A��.��=�R���u��������ƻ�:°�r�����P���鸵����R��������R �ϾI�I ��Iђ�TVSP��� 3ҋ�S�<�6. �<[�<���6. ��;[^�T3ҹ @@��V2�ô ����������<u2��0�@ �J���\�L�6���$6���<�t��2�R_���te�u�*�A�  � r\�� u4���@�*6;\htɋ�3۸ �/<�u�u��/���/
�t��ð���6�\h��� �����\���,�� ��s�<�t�&����< ri��u��
��1< u���FE���D�$<#u"3�.:�Gt.:�Gt.:�Gt	.:�Gt@@룋�<!u�t���
E�D�����<"uE�
�t���D�D����rx�*���u�Th���u�\j;ThuQ;\juL�\HQ�LJ�v:t����Y��x��Y<t� � �ȋ�����L끃�9s�&������� ��2�P]� �/<�t�빸�/< u�DH�����*<u�\j�TH���\�T�<u3�Th� �/<�u'��/
�t�<Au�A �$�&�'�#���뭰�����^r���r�2��B��T�L�\����������6�,6�.�!��\�L�6�,6�.�6�6Ê���� ^r6�66�G ��1 &�����\�D��! �&�&�_�6�� u�6�>�  u6�� �3ێÊ������
��/t<��t����T��$�>(�&�.#���|
�D�\�L���V�*6�Dj^�
�u�q��D�.��=�D���AV�Y��Dò ���]r�r��&���2��9��L�\�|�T����&��D!�T����D& �Tò ���B]r"�>�&�ED�u��8I��r���l�D2�ð�ð����L�&���  ����  � ����P� �/X� �������| u&�E �w�Ь�Ȫ��2�u�������Ī�إ���������H�3����GG��&�F����2���&F��&�F��&�~ u2�\�T
+؃� �t����������&+F����@��&�F&�f���r��u��=�r��҃�s
.�6�MH;�v��&�F&�F  &�F���.��=����0V�
���\�6 ��3����� � � �64 �.��=�>� tM.��=3۹ �W��r$&�Eu&�e�����pt�>����	�UW&�&�GC�̋0&� �0��.��=�� X3Ɏَ¾� �
 � �&� +�=�v��- � +ر���ڣ � =��t� � �   �  � � ��P �!�R ��4  �6 �2  �8 ���: ��&�@ ùf< t<u	�F��qð�#�VWP��4@�@��&�G�(@�z@:�u
�u�X_^�P��@�f@�
�u�X�P��
�u�X�WP���2����X_�� ���� ����6�>r u�Q6� �Q3���Y��Y�U��S�^.�8^s�^2���C^.��^[]���[]� .��=&�>����t&�ED�u���&�E��.��=�2K�������&�E��;�t�t�����t��&�M&�5�:�&�����ˊ��7^�6�6�6�6�� ���W6��6���6�j6����6��þ(.��=�4�D"�\$�6�6�6�6�������6��6���6�$�Ü6�> t�����P���*X������Ü6�> t�����P���*X������Ü6�> t�����P���*X������Ü6�> t�����P���*X�������V�x?u;6�>�
 u��E2���*6�>��uPSQR�  ����� ��ZY[X6����2��2^6�� < u6��Ë�<$t������Ў���2�
�t�܊�:�v�8t�݊�J6��6��V��6�.y�����c�<
u�\�<t�.:�GtC<t6<t2<��<��<t2<
tD.:�Gtk:�s�����6�>y u�:�s�F����a��A��q���8_�u����������J�
�t��; ���6 
�t&�E�<0r<9v� <ar<zv��h��\��^�6���\�9�� �O�
�t�X &�< s<	t<t<t�E 6�>y u�
�t���N�WO��ΰ S���v	&�}	t	����6*�*�ˀ��[_t�� �����O��x� �s��n.��G����*���4 ��6�y :�t:�t������������:�t���F��� �������.:�Gu������*�tItW��G�_u���*��]�j��@�� _W��^�����6�y�N���v���� �
�� ��<�t�C�6�>�3��T!r����/u��<&�M@2��&�e��<S3��2![r��/u���*��2��/�S� �!r�\�　��� u�\�Gt�)�[�� ���� r�P��l<6� ��;��g/t�@Xt��\/��VW=  t�l�Z��l�Z�Ў؎�� �_^����P� XÊ�< r\<t6��V6� 6�& ?uP�,<X�X�^6���t�SV� �a r!�\�ǀu�Àt� �L r�Dt	6�� � � <t <t'<	u�6�����Q�ȵ �� ����Y�6�� ��q�6���v�< s�<	t�<t<t	P�^�S�X@�M���;� ��r���Z;��_.t�2��X.�S� �S� ��P�k;XV���^[��^;� t���PR3��r��%.ZX��<t<t<t<t<
t� ���c�� ���D!�T#�|@s�t$����Ur	��r���������V��T^r�V��^r�Ӌǋ\�u�� ����3���P�����Z� �� �D!�T#
�t��t$�2��t�D�6�k��r�&�E2�P��\u6�k&�E�D&�E�D&�E�D&�E�D&�E&�M @�X�>�Y&�M�&�= uP�M�X�s�<t�����R����>�4V����'T^�Zr6�6�6�6����Tr�r�����6�>��S�t&�E�D���g�3\t�[&�E�uB&�E�D&�E&�]������
߀��
ÈD&�E�D&�E�D� &�E$�&
E�D
�t*�&�E�D&�E	�D�@��6�� �E�6+@ S�;��D[&�E$?
ÈD6� @&�Eu� � 6� ø �W6�>@ &�M�}&)w&���;��_&���Z�.��=
�u�>]>_t�>]�>����� �>@ &�M�}�����Ӌ�&� tN&�=�tH&�E �u2�'[u-�>]�_
�t�&9]s&�]����;�ʋ����u�����u0�Q&9Us�&�U����
�t���9>]u9_t�w�3��]�_�l�
�u�>]�_�>���&�= t�]s�<t���2���j�.��=&�>�rð#ì�7���ÊD��t�yZu	� �/
�t6�:��t����]Zu�P� ���Xr�&�E�$?� @�L����
ŀ�&�M&�E6�<&�E1VW�K� F���k��'_^r&�}&�E 6�6�&�u&�]	��&�E%? V�NP&�u&�]	^r�D&�E�D$�������
�$?&�E�D$?*�&�E�D&�E&�E5�D&�E&��t�} � ����W�; �_+�&�&�EH&�E��D�tP6�>@ &8ErE�;��}�6�<&9E1u2&�= t,�D��t1P$�<�Xu6�� r�&;]u$?&�e��?:�u��ËD&;Eu�è@u �\&;]u�\&;]	u���PS�D�~�[X6�>�6��s����`���6�$r�6�>�6�6<&�E1�.��=�# &�K&�.�� ��&�V�8�ËD!�T#��@r2�ÊD �T�����؊��2��PR��$�D �����ҊŊ�DZXË�<�u��;�Ë\�u��� �\�U����F��F� ����F�u� �N�������^��F�t�|��F��V����F�����F���׉F�V��F���F�6,�� t�F�6�,��uH3���F���F�3ۉ^�9^�u�F�t�v���s�U��F�  �F��� �D&�E�D&�E�F�V�&�E&�UR�N��q�F�u�,tUV��^]r�6�> t
6� �F��N���&�E&�E�D&�E�D�F�3��v��F�F��V� ;F�t�F�u&�E�u�F��t&�F��V� �F�t�F��F��N�+�2�6�>,~��V��F��F�t�F�t�f��F�t�D!�T#�|@s�t$�F�u���D�T�F�t	�N����L�F���]ø �`jRQP���[NXYZs�+��(�P���Xr*&�E �VS����[^6�>�sP�R���X= t=$ uP��X���i�u�TVu
6�>]6�_&����&�E�u	��tM����D� &�E�D&�E�D&�E�D&�E�D3��D6�>@ &�e:DtP��Xs	��:�u�2�ÈD&�6� &�E�>�&��V�C�?��ܹ4i3��W�t�D����
�e���`���[�� �V���Q���L�6��6����<�u���4���:Ms[���6,�6.�,��.��.�,s[�پ��>��l�t��[
�u�6�ì��G�
 �ê�>,�l�t������ �m��ê� ���6��6��6�m 6�l ����<�u���6�m6�l�P�D��
 ��6,�6.�,��.�c�.�,r�V��>��l�t��[&��*��6�m���Ls�� ��6,�6.�,��.� �.�,s�ھ��>,� �V�D�����FF��^�5 ����6�6,� ��6,�6.�,��.���.�,s�뫹 �&�}� uOA��r�<  u�| t�.�� �&�}� uO��3���6� �������Js��.��=��0�V.��=�6��DC �u .��=�L ����!W^_ră� tO�<\uFP�
�t<t��<\u��<u��
�u�X2��4����R��W�qK_sZ��6�>z�u2���Jr��t����Z���Z�q� �����,Ks���>z�u��>����t��Tr��>�&�EC  t%WQ���|�\����2�W��J^�>�&�EI��Y_�R w�&�EC �u&�EC  t���&�MI�>��,�2����o��V���J^s���6�>z�u�V� ^v�����r���6�6�Q���CY�\a\a�a�acc�a�ahb�b�b�a�ab�c�c�ab��<wP����� ��X.��a��+Es���< &�Et
�t���t߀ʀ�#&�U�h��#2䨀t�#&�}&�e������T����Dr�&�E�t��#&�}2��K�,t�P�Xs��:"���u���Ɖ �tu� ���Dro&�E�uc�#&�}��#��uN�uI&�E@tB�~<|&�E�t2�~W�|�}�.����6��>����6��|^�� �������1u�&�Et�6�~���6�|3�6����|V�W#^6�% �	���K���HrH� rC&�U��6�>�&�ED�t� ����A��D: � ��*s�� &�EDt�� ��߉T뮰� ��Cs�_�&�U���U�� u�&�E@t��~�t�~���|3���������6����|�"6���u6���6�>��� ���k16�$�P���HGr$2��#�>�&�ED�&�}Eu�#&�]&�}�X����rW�>�&�ED�_�X�B�������u�&�E@t��~<t�~���|3�����|V�"^6���u�6�}����u�s��/��o �*��~ �6��
�u����<*.u�|*t��	���??� �u���=.?u�=??u�m$<u� �L�su
�t� ����ø ��u�> t� ��
�x��o�&�>�6�ku	�Gt�2� s�*�E@u�6�M@�'��o��r&;^w�)rS�� �.��rG�4s��.�&�F �A5r5�ot'�ktPW�>�&�%��A�&�
2����1_X�7���ou�=��P�WPSV6�>���6���߃����I��/HG6�>��^[SV�� ����e2��p%�>�&�E &� �5Nr�>�&�  �"N��.�^[X_ÜVSP6�6���2�X[^�ÜVWSP6�6��K��2�X[_^�ÜVSP��Ծ26����s��/��#�6��>���%  :�t� ���6.�6,�.�, �p ���s= u� ��,�.�"�ø �6,���Dt�6����w؀>p uы�����s�  ��V�6,���Dt^�^� ����6��6��������~����r#
�y3� ��P�v�3X�>J u��s�X� �k�u�>J u
�u� ��X��W�K� ���d�5�K�W� ��k�~��Bs��d�.��r��s��>J u*�d;/t]�@�u�k���e�6��D 3��"s�T�S�>��`L[�>�&�E@u��3&�M@�����@� ��} rw��������m rg�����K� �>�&�E@u�3&�M@V�6,���Dt���^�^�!�r��~ �r!�w�Y�s�  ����@�t���������������/�.��r	� �-��ì<?u��C����X�s��/����L�� su
�t� ���ø ��
�x�>��u2��������3ۋ��L�T2�D�u�|�\������t�#�'�&� �����sP��/[���P�L��s[�
�yX����X�>��t
�j�s�  �:� ��4�>�&�g�&G&�E@u�V2&�M@�vRW� �Ћ����_Z�21s� �O��6�:�g�6�&:���.��=&�>��c�u�9&��2䨀u�t�� � �Pt
� �#�g�>��6����u��tP�.�/[�� �P��/[�&�DC �t� r&�M��u�P��/[�� r&�M���rs��
����i.��� RP ����m�t�>�&�%��A�&�
�� �N���,�h� �>��� �Z��P��.�PW�Ċܰ�f�lSR2��$�Z[r$
�t�K�������� �F�2����_X�6��tP6�&	EX���L �@r+�>�2�&�E�6����u0��t�P�.�/[�� ��� t	�t�#P��/[�&�DC �t	��u����w�:�s u
�t� 6�&:���z�� � �� ��t�
�x?��&�G�u�t/V�6��L�� �u
�р����pu����L����� t^�^�6�&:��J s���$� �>��� ���>��&�E �t�0&�E1�&�E �u&�M����� u�Hs�  ���� Q��GYs�����>����s���ânS�؀���>r�u��pt��@w�؀���w[�ø [����s��/��#�R���*rA� �)r9�6��d&�N&�V���t;�r#3�I��(ruBC��KK&�F��&�N&�V��)�Ë����>����u��/�&�EC �t��/����� t�:�L�Ds�&:��su
�t� 6�&:�����ø ��
�y
�H���p�>,�6��,@��>,G�:t�����K�&�}�u&�E��
 ��k�P�H������X
�x�>��u�:u	&�E����|�����  ����&�=u&��6�&:���4���>,&���t��/��#��������@�<r6�>�&�mE��&�F �v�~ ��L�6,��K� �6�k��y���P����.��sX���X�Dr��sr�2����6�6��
�t<?u���6�0&�2 ��QK�Y9Y����/�� 6�>@ &�M��}6�<&9E1u&�  ��;��3�S�8[s�&�=�u6�<&9E1u6�>&9E/u&�  C���>�&�]�� �t��/�����p�� PS�dE[XP��� t� �� �s� WV�t �����^_t����� �D �t&�m�D6�k��D&�E&�M &�E6���D&�E�D&�E�D&�E�D&�E�D&�E&�G@u�f,&�O@V�L6�vR� ���u��|�L�t�6;�t�6����Z�+_�r���P�Y�Iu&��-�Ü&�HuH&����#W&�U�&�U�6R�\'Z�r%2��K��)r^6�>�&�M�ߍ}� �d��_��>�&�]��� u��� �t��/������ �������������� u��� @u�PS��&�E&�U3��� [X���s��/ø ��n���j�����D����>�q  ��r�= t��.��>�+�V�u�u�6�3����'rw�rr�>�&�E@u��*&�M@���. ����..Z��.��KZ�2���(rc���>��M^��3҉T�T�E@u�*�M@&�F �)� ���ZZ��.��K2��y(r�>��M^���������^����s��/��R�&�EC  t&�EI���L �m�:�t��&:��� ru;����<���S�s��/����L �m�Bru�>��u�	� ��XXX���>�+�S�u�u�K�?� �2����lrԎ���=. uȃ��=..u��H �Jr��k�=s��>J u��.�����r�Z��K2��n'r��>��M[���������W ��WP��������X��>�&�E$<u�"����x�t��/���&�E�u�#����%���#&�]�>,��@t��t2��� �� u��ta�6�0t��t� ��3�����6�6��g�״�6�>]�y#� ��6>l6+l
�t<t��_6�>��{_��6>l뒌��؋�3ҋ�Q� �Y6�6��t��W��6�>]�y�_6�l <t�<t�2��_6�>lu6�j�6�h6�]  G<t<�@� ��3����5&�G6�6��&�G �t���T��
�t_<tI��&�G uG&�G&�G 6�6��p�״�&��� �t���
�t%<t���I�&�G�_6�>��P���*X�~�6>l����<u�
<
��u3����	��6" �>�u	�>�&�e��������6" �u��>{�t�{��QW�{��_Y�}�<u���O�
���3���>�&�E$< u��&�E�t&�Eu���=�t�	�/�&�E�up�#����r�>�&�E@tQ�
�Y����3��6�6��[�״�6�>]�y �6+l��6l��
�t<t��X���X�l�>����Ë�� �#&�M@&�]3������,��3Ҩ t뎨un�uЋ?t�Q� �Y6�6��t�k��W��6�>]�y�~_6�l <t�
�t�p�_6�>l tB6�hG6�j�=t	6�]  ⳋ��\��~���Q�<t�t���X+��c��>�6�>W uW��0r�Ǝދ�_Ã�w�6�6���3҃>� u����&"V&�N��s�Ȋ�����Ԁ� � ������%r����s����׊���K2��+#r�V�6��L^�6�K��&�N&�F2�R6�  QP���] XYt ���Z���O t�6�u � <t�<�u��Z�&�Et���Q�uI����<Ys�gs��&�Et��2��<s�)s��Q&�f&�FS���'� t6�u�: <t�<�u��Q&�f&�FS����>�v���[6�l_+���6�]� ��<uP6�p6�(6�r6�*X���&�u6���6��,���t &�E&�U����&�E��u<�.�&�^ �v&�^Q�A�������ы�&"^�s�NYu&;Fw����,s�,��uH����3�[�á����t&+F��+�s�3ۣ���3�&�v������u &�E�uQ&�M����� Yu�|;s�3ɸ! ���u��&�E&�]+��r&u
�t ;�s���t�s��.��~�����r�t��%� Y[3ɸ �É����>� t�r�>� tS�r��t�s������r�WPS�K8�.RQ�"���YZ6�r�6��^ Y[��_s%� ���á��t���Sr��  �s�l��>���+,&�E�u��&�E5��&�E�	&M&�U ��6�>q  t<6���ʃ� ���E6��&�F :Eu;]u;Uw
;uu;Mw
6;>��=u��P�E@t/QRVW��+E�؍u&�N��6�>�6����� �_^ZY���t6;�Xu�����s���&�e��&�E�&�E��.������������� &�^������R��u- �� ��ZPR�������ȋ��t �� ��3�����X�>;>rgt+�>�	�  +�rVtG�ʓ&�f����&�f�С+��� Ã� �$������s��v3��>����F�� +�v	3ң���X���r����+�t �Q���@Yr���BIt�{r����>� t	����r����tp��� �Ar_�t�s�����\rIWP�-6�.6�K8���t<'t#6�u���<t�<�u�Y[r�� ���Y[���'������t����r���  �cr��>������u�&E&M� �� �a����tk- �� S&�^�[�щ�8���jr��&�:r�>���&�E��&�E� �� 3��4����>�&;Us&�E  &�U&�U5����r��3��>�&�]&�]5&�]�tUPQR�.�&�V �˴���ZYX]�|r��SQ6���ʃ� &�F 6�>w  t16:�u*P6��6�>�;�u;�v6w �� ;�u;�s6��  X�v:Eu';]u;Uw;uu;Mv�E@t���E� �^��=6;>�u�Y[Á� u�ʋЁ���Ċ��2�����Ëȋ�3������&�N2����������Z�k$�<u�~�s� ���'
�t:6:&t3�Gt6�{�֎Ƌ�K6�>K�u6�K�a t(�.��f s��P�H;�s��:&t�����4�,�&k�䞍t��t	��t�2����t���t�~�t��.�&�f ù �t&�}�?t�áH;�t$@�_ ;�u�s��:wr���Ns��r�2�ãH�Ès�H�>��U6��U��6� �"�3��$�H�H�����%����&�^������S��[r������&V���t<��&�F���wV�:u��s^É>���2ۈs�P^R���Z����3����sH��&�F&�V+¢w����  ���~ ��#�����>��}:\t:����� r.�m�k�#�K�>��׹ ��< t������� ��������6����u�u�k�>����&�]I�6�;�t@;�t<�:tBWQ�t�VS�D� �6��0�F�;��_r�< t���[^�D�Y_s�6��t�.��?�.����r�E2��Ë��׎ǿK�	 �<.t��t
�t����Ã�� �Ў��������< u	�m�k2��V�����>��t;>�u�>�&�MI�Ў��K�  �������K2����<.t
�t$<\t <?u�����S�
�t<\t
<?u�����N�̀ɀ_;�u�� V�
�u�>m�>k�0r
�t�� ^�|��>K�u�KWQ�s��Y_s�� �>��Gu� 6�>L t&�׌�_�:t�:t�>f�= u� W���ً�:t�ڋ>�P��X���=+�+�SPVQ�u�u���e��Zr
�K2��tY^X[s_���!�=��>���_��
�t4G���~u��N2��,_�:t�:t�>f�
�t����h���^���
��m�k���.�3��H�{H�����P6�k��"�$X�VWQP�6K�>Ku�K��ku"�H �D �t�ƃ�
�K� ��t�4���u���юُKXY_^�6���|������6�6��޸  �S���@�3��
 ��ǿa��������������K2��U����~�6�6��v��^��M��DC �t� 2�6�L�΋v��,�L�>�U�]rn�6��|I�uV6�6�;v�u�~�6�>�����6mU��][���m�v�s6�6�6��3ɈL�DI��6�6��DC  t����LI�~�6�>�6�������~���]�WV�����uF�  =deu-� <vu&��u V���< �u�m�k�|�^_s��_�����6�:u� 6�:u��06�6��F�;��_rg�\�6;�t]�< uQ6�k6�.m6�.k&�m��YuO6�6f�ًG6�H�G	6���G6��6��&�'6��  6���ߍu6�:�=��u6�: 6�&:��Ü6�:ty6�:t6�&:�6�>f�^SVWQP6�>��;�E6�D�E�D���D�H�D���D	�Ã�+Ǳ �������} tV[��0&�\�XY_^[6�:������
��6��6���6�� 6���D�t� �D�u� �#��ڌӎێ�3ۀ�u�� �3ۈ���.�����.����|�&|�.~���o6�>#�x4�Ў؀�u�����&��Ԁ�譽�6�� �=��u6�� ��6���Ê���<u舽�K�6�&��<u6�� �
�t#��t��t��t�t� �D�D��' �0��U �� 6�@���6�&���= 6��u��6�l�:�6�6,6�6.6���6����.���,����l�.�,��6�&l������&�E�ug2�&�E�&�}u6�>vR&�e&�&�}&�Et@���Z��P��X�આ�&�  P�) &�#�y�D�t��������<uX��X�d���t���D�uM&�t&�t&�	u8� rU�Dt&�6�n6�n��6�t6�6�v�6�> t&�G��"�D6�x6�z6�x�D6�x6�x�Br��2��WQP���Z�X�P���3����X�આ�P�ë�ثYX������_�Z�WQP�6���6�>w  t!6�>luQRVW6�n6�>\t�� � ���'r
6�] ��k6�6�n6+�6�=  uR��wM6����6�w 6�l6�j6�6�h6�6�s 6�h6�u 6�j6��6��6��6�n6��6�6���6�6��6�n6����_^ZY�6��6:�u6���6+�6�=  u
6;w s�������r� ����6!��6�>� tN6�6�j6�6�h6�� 6�l 6�^�uVWRQ3��1 YZ_^�6�l 6��  6��������g�rA� ��6��t5��6�&�6s 6u �ڋ�6�j6�>h6����6�>j  t��f����á�=��t�Ã>� u�Ë��t�^r� �^r���u��r��H���+S���p[r��QPU�&�V �����+�]XY��2���&�N��2�Q�K���wsY�&�N�>�&�MW��3����s�_&�E@u�W&�M@Y��� ⺡H@�ë� �  󫪰���
�6��D��D��«3�����~��P�L �m�K��ы�Xs.u���t�2�����t�����u�� ��>�3���ZtH��ku;
�x
�u�Q��&�o��u$��Yu2�2�PQ���F�>�VS�*sZ[^YX��Y�둰�P���t Xs������r��ku�PSV��)^[Xs�P�>�&��&�E@u�Q&�M@�.�&�F �5X��>�3��.�&�PW��)�_&��;�[^YX��r�PSV��)�^[X��.�s�>J �u�� �r���r����
�y� �-r��kt�>{ u�����K� 󥤠k��3���H�����3�W����6�&�D@u�&�L@�.�&�F PSW�>�&�E�uS��&�]��&�]	[����
_�\�� [X^��sÊ��>���2�
�x���G�3���@��G
�x6������V��������ȭ
�y3��ȑ���3���
�xD��GW��&�E5_�:t�;�D��D����6�6��D��D��Ã�+Ʊ ������� �^���>���U6��U��r5&;Nw/+�S�6R����Z�s[��K2��r[r��C�������P��>�
 t��
 W�>���_�X��>�&�]5&�U�t$+�s�3�&�]���r������s��B����AJ�Ë��s�K8�Z��r��t�6�������>��>�&�M�}>���3���s�-�Î.�ۇ����� �6�>��]+��W&;vr6�>m �á� ���� ��;��wr��;��w2��]�r��.���� �6���G@u�T�O@�w+�&;~r6�m ���t�t&�s��&:Fv����s��r�>���� �s����RS&�F����*ѹ  ��r7Ȁ� ;�s3��C;�t�K��+�R��&�f�6�ƣ�XZ+��[� ���Ã���+�*��̈&s����Q&�NJJ6�  
�t2����6���
�&V6� Y�6�6	�����s� S3��8�>�[r�QS��&�^��w	&�F � C&;^w^�r/u�&�^�� �Vr &�~�t&�N��ڋ��Ar����˺���4[Yr���r��9 r����t�R&�V �>�&�]&�]5Z�&�~u�[���� X+�� ���SRW3ۋ���_Z[�3��r$t"��R��Zr�u&�~�t&�F��Ht�Kr�&�F VQU�y]Y^��Mr�S���.[s����6�N 2Ҩu&� G� ��� t�3����t�3�󪑫�����t	� �(uF� �� v�<:uF,@vP�tXs
6�>t���FONG� �( �<.uF6�t�� �� � ��6�&����N�� v�N� u6�N�t< u��I<*u�?�<?u߀��ڰ �Nì� t�N�6�N�KW�  � ��2��Ъ_�z�6�>K�u�6�K�fffffffffffffff�����O�n�����DD��������������of�����������������S�1<ar<zw, <�r
,�.��=�P� �X[�S��P� �X�P� �X�<~sS�ҏ��.�[s��������$ð�</v<\ð\�t���  �    6�>!t�QSV�ӎÎ�6��6��6��  ��6�62 �;�6��t2�^[Y�6��<u�6��6��6��6��  6�� ��^[Y�� <u	6�>� t�<t�� �6�>X t#6�>  u6�6X6�> u�(�.�|�6�X���F�S3��C�[r����t�<u�6�>� u�2����J6��S� ��[r�W��&�EtP�&�/Xs6�� P�$�/X�6�>� u�������_��b���g�t�S3����[r�2��W�<t�<u�6�u����>��>W t������&��`�.��=�! �  �&2�2�> u��#��.�t��P��.��=�
X�:�X;&2u
�:�
齮���t�
� L.��=�M���xG.��G.��=��� ��������  �����6����62 �W�&���&�� �6�>  u��6���u��86�&K6��6�.�V��� ���d ^×��� �� u
P&�F 6�"X+��R&�fZ�2�&;Vr��&;Vs&�F���
��&;Vr����6
&u6
&K&�F 6��6�.�&�v�����v� 6�>  t��l6�&�6�>��tV6�6���^�6� 6�!6��t��)6��&�&�&�> u�$�.�x�&�&�&���Ŏ�6�&�6�!6�  �6�.�<r>tF<uL6�KtD�6��u6�J6�"�6�>��u�VP6��6�6��X^�6�K t���6�Kt����>W t��݀>Y u��|2�����*6�Y��"�/�"�B�YS6�0�ۡ ;�t;�uP6�>|t��U�6�0���¼��ܼ�U���! �"��Y �����0�0 �&. 褭P��.��=�
X��XXX���$��P�6��6����
�P��-�.��=;���s���2�$XV�[�<�^�&�~�s���t���Ã����u�>� ��&;^w&�� r�=u&�v���r�������������&�F��P��6�K�����<�u�X��u�� �� rҋ5tQ���Y���&�~�s
�� �����3��56�6��D@u��L@6�>x t�PSQ�������$P������ 2��]Xr�>��E@u�U�M@��O&~��Y[X��x PSQR��&�~�s��3���&�N�� u�Ё��������2������&FIPRQ���  2�� ��YXZrW�6��|�;�u7��x������  B�  2�� �r$�6��|�����ZY[3�&�~�s�èX�ZY[X�&�m&�F �v�'��y �W&�mE&�F �v���e _r�u83�H�G 2�&�uE6�>< &�ED�u&;uEu��&;]Gu
&�EIt&�EI��X���.���&�F����� �K��v����.�<u���&�f�Z�\�]  &�F�g�Z&�v���>]�x�2�&�f�v8�
u��
�� 
&hy�et<��U&�n&�F]t&W�K�>i�*�>(� �u��_<t�n�6�>q  t�� 8Eu�E@t���Ë=69>�u�&�F���� 8Eu�E@u��E� �� ��=6;>�u�6�>w  t6:�u6���&�~�E u� ���r��>��U3�6��z �E]r��6�j�>h�&�f�Z�\�]  &�F�g&�v&�v�Z^�R��>]�x)&�F�6l&�F  ��6�>h&�F�E�&�F�E�2���J�6�>m 6� ��6�>���5� _�PSV�6�m ;�t ;�u6�m ��u���D�w�<��u�^[X�}�u6�>m �;�u
QR�ٌ�;�ZY�3���&�F �> 6����t;Uu;Mu:Eu� �o�;Uu;Mu:Eu� �=6;>�u�QVRU�]Z^6�s� �2�68&�uJ�]� VWR6�>y  tS6�z �t�[ܴ��ܴ �6�>y  t&�N�靋�_����Z_^rH6��M�U�m�E&�F �E�E
3��t&�F�E
&�F�E���6��6�  6�>�6�> ����6�u6�>q  t#�, �e68&"t6�t�E� �=6;>�u��>J u��ô�8et�:�t:E�u��E@t�P�u� Xr�俉EXø� �E<�t���@t�� 6:"t�6���m�]�U�M6��M
2�6�K��t6�K �EW3�SWQP� SR6�>y  tQ��&�N��6�>z ����Y��Z[XY_rG���[�u�_�P&�F6��&�F 6��X�6�q �6�>q  t6�q �3�6�4钨6��  <uY�BQU���<v6�#���]�t��T�<t�<t�<t�^��F��F��F� �V�^���o��N�6�6�� 2�U6�� �I�6�&� ��]r��F���2��f�r�t
��� �
�� �F�  �F�  �F�uT�v���u6�0�, �t?��3�� �2��u�IxƮu�W�]^����ZYs�t���F�3���� ��v�N��� ���rP�tL= u����u�F����=MZt=ZMt�������+��F��F�tI�~�&��F�&�E�F��� ����^��D蝴PU�i
]X��6�6�� 6���@uԨ@t�6�� �)�F� �>� u�>� u�F�=�s ��t�@�� ����w��  ��r�;�w��F��u�r�;�w�+��r;�v���؉^��>s�q��� ��~� t�� s���� ���F� �F��t	F�+F�- �F��F�V�V��R���X���ȋ^�2���
s����^�� r��)^�S�����^�3�Q�YrH;�[t+ȁ� s;^��F���uŋN�������������������3ɋ��^�3��
s����R�����Zr�c ���v��t&���F��7��J����PQ�F�6��6��6�6�bYX�� �1��F�t-�v���F����c6�6�� 6���@uب@tԋF�3��z�6��t6�@������tǉ^�S�[�F� �F�3��� s�ñ��= v�- - P�^�3ɋ�3��	Y�^�3�Q��^s��;�u�y�6�� 6��F�u2�F�- 6��6�� ��� ���t�� 6�6�6�����  6�a �^��U��]��F�t:����6�>? t&V6�6@&�< t6�06�6�&�@ �6�? ^��]�K��V� �F��tH�؉�F�H�؉� �nQV�<.t���s��2���s�^Y�iR�v��踮Z�v�&�, 6�6�&�@ �v�V�t� Q�\ ��3���Y^V�t
�<󤫫^�t�ɀ����Ɋ�2��e
s����2��Z
s���6��t�t�t�t&�
 &� 3��؏� �� 6�,� 6�06�.�F�t'6�6��~�&�]NN�&�u6��&�]&�E��]�E�6�6�6�>���6�> t.��=�� �c ��P�P����6�! �Ћ��V�ڋ��� �^�U�A]� �S+��6�� [�S6�0� �E�[ÜP�F��	 �F�� X���t�H�؉ ��v�ά<:t�<\t�< u�+���I6��6�>] ���t:&�
�t36�>:�uGQVP���u��X&�6��^Y�X^Y6�>2�������P6�|6�0��s� ��S�9[r��ã X�&� 1���ڱ���%�2�6�&M
�6�| t6�|蕠6�60�D�2�6�| 6�&|6�4�w��\3����
 �� ���������6�$ �  �0 r=9 u�> �=Zt� ��6�� =��t��;�s�ь� @��&�=Mt&�=Zt�À=Zt����r�&9> u�&� A &����詮6�$ 6�� 6��t6�� t6�� 6�� 3���6�@6�B6�DP6�� ��r69> ti6�� t6��t6�� 6;$ u	��6;� ��=Zt�V�s�X�U����6�>@ t� 6�$ 6;� t6�@u6�� ��Q�[�\�"�����-�r�� Z;�v��R;�w�6�>@ u6�@6�>B t6�B&9 v6�B6�D�R�6�D� +ˌ�tLю�I���.3�6���?���w�6�@r6�B� +ˌ؋�t�@��I� &� �M�&�&�> ��6�0� ��@[�n����H��  ��H�a�s�����g�r�� Q;�v����$�6�� t6�>�  u6�� �  ��H�'�r
&�> ������	鱟
�t <t$<t2<t66�#���6�#���6�2���S��?���[w�6���6�� $��6�� ���t���rt�6�� t�) r��  Z6�&� ���6�� u� r��  M6�� ��P6�$ ��3�&�=Zt���k�r(6�� u&�=Z�;�u�6�� u���J�r;�u�X��X��m�֥n����������;�;�;�I�<r<	v��\6�0u6�>�\6�<.�6�.�6�P��6�#�鍞�3��ūS�+r#&�= t&�=�t&�E �u�>������[C��蹫[�L�6�� r���6�� ��6�� ��6�� r�躜�\�|
�D�L��XV覜_�H�V� �GG��^��\�L�T�|
�D�t�\^6��6��6�r��Y�� ��
�:+�+���� ���R��D�|�T�P�%�/[r�鱝�6�$�D
6�(�D6�*�D6�&�D6�&#�.��=&�0&;2 r���&�>4 �����r�&�=�u���S&�2�� [�.��=&�>* &;]r&+]&�=���u���P�; ���X���3���r	&�=�tC���P3�S��[r;&�= t&�=�tC��6�>&9E/u�6�<&9E1u�&���6�>&�E/6�<&�E1X��X���[r+�>���&�=t
&�E$�<pt� �&�����r�>閜霜�(r�>�����r�h����3��s� 6�0&�2 ;�tPw"� &�6 ��+ˀ<�u?F����w	� � S����t}�S����ہ��U���]rd��3�6�0�� t
YQ�
뒰됋2 ���64 �YQ+ʰ��6�0�>4  uU�6 ��]�� t�4  ��4   �6 �2 �[�뮰����q�-�r&��As��6�>�6��&�E t6��6�6,6�6.� �֏.�,s�ʋ�뫋�Q���Y��Î؃�6�,6�.þ,t��� s�<v
6�#��<r
w&U&M���&�E&�U謙�T�&�E�u
&U&M��&�E�u�&�E%� =@ t=0 u޸!�/s��<s@�u r�
�u�&�M&�U��[��L�T� ��&�M&�U3�6�� &�e�&�M @���6�#�밋��o�rW^�� r蹿���&������SQ����[X��������rP6�0t3��6�>&;E/Xuð��<u&P���^Xr�|E t<u�LC @��dC���� �<t�P��/[r����6�6& ���t	:t�t����P6�>�&�EC  ,@68F r6HPA�:&�&�E\ &�MD@+�&�EI&�EK�&�EOXV��r&�uE&�]G^X�P,Xrt-<v<6�#����6� ���L�� �3���r�6� ���6���P��/Zs����� r�V6�6��DC  ^t�6���
�u6�6@HV6�#6�r�t!PW6���6��A��&�EC @_Xt�� r�DC @u�6�6�#�^�6:G r��SP6�6< �X���6�6�6��X[��U���W�~�6�l 6�m 软t�D�6�m6�l���V�r*�z� V����t��^����_�v��? tU� ]s����]�2����6�L��6�q6�z�6�>�6������� 6�r�t5����r*��]�8r��6��q�t�6�>��E�����_���6�����#�/s)�P��R���M�u:�uX�����
�t�:�ߪu��� ê��X�< u���PU�  ]Xs6�r��e�6�r ��/�蓣���'��/��r�VW�[�_^�r�V6�6���\O��� �r�O�\&8E�t�O^�� u
�t�����t�N
�t�\��S r��>��6��u�D���t&�= tG6�>��6�3��q�t�,�>�&�EC �u��1����K��ì�Q�u;�s���N3�8u&�}�:u�\��Ī�����t����Q r�&�=.t&�=..u
O�+ �r���� uҬ� �u�;�sȪ����t�N멊
�t�����;�rO&����u��ð�Ã�VWU��.��:�u���t��:�uW���uR2���v�G�v���;vt?6�r�u��6 z-u
�t/�v�K�~
W耱_��IN;N s���~������� �u��]_^�����I��6�Z �tj6�6�6�6�V_3����rK���DC  t�W� t_��&�= u6�L�u��_� 6���x�+�6���< u�\�膡�����6��6��3�6�6��|E6�>�6���VWQ��������Y_^s�7����=��#�2��< tӀ|:uͭ ,`uư����@�:���/�I�u�P�D��k�t&��u�Xì�o�u��X��2��]�`jP������6�r6��6�>�6����s� 6�>�6��6��6��&���Q�<�[6�6�r
6�>z�t��PX3ɉL�L3��`ju	��t$� WV_躺_Q��Y�6�r� 	L6��6�� 6�����7�=W u�[�  6�6�����Y6����6�>$%u����Q�4i6�m�'���PQ����YXr3�>z�u*�m,rt�#������r�[��D닋��J�r�����Q���[�Yr�6�>z�u�� 観r�ذ��QR���>�1�6�6�6��^Yr�6�>z�u�Q����Yr��>z�r��6��6���2��k�r�*�t�������6��6���� ��r��Q�j�����P$A�X��u��U���
����t� �m�N��V��^��^��������u���3��O&�E��E�t�\��~�U�ȗ]�~���������2���V��N�U��]s<Pt�<u6�>$At
6�>$St�����]r递醒6�r�u��6�m�6��6��  �� �uE��� t>����w6�����w.6��6�>�6�6�6��6��6�6�6�6�֋����Y^������  t6��6��6�&�� 6�>�u���r�6�>� t
6�� � �Б6�� u'��r�6�>� t�6�� 6��u[6�� �R��6�r�t����s26�>� t�= u�6�� u�^6��6�6���`�rM6�� �6�>� t6�� P�ݏ6���DX��?�[P6�>�u6�6��s���`�X�� �� �!�<wW��s_���6�#���ؽ��V �NY�N�v� �ըu�&�E�t�
�/��� s�ɡ�Ð&�E�t�
�/���� �� SP�� X[s�ݜKu���WQ�! �K�.�� ��&�V�b�Y_<t���.��=�> ��� �W�u �K�.�� ��&�V�)�_<t����� �Q� �>�3�&�E3Q��Ys
�\�����s�YË��D t�D ���L
�D6�6�b�D uV�t�,��=�^�D6��&�@ 6�> t �D6�� �D u����6�� 6�c 3����!`3��C���73��� �"��fPQ ���YfX�X�̸��g����X��.f�  .f�6  ��.f�  .f�6  ���RQ��f&�YZ[�fPfSfQfRfZfYf[fX[`�  ��af`fa�Z� ]�   l� p�	 � �� �� � �� �� � &�>  �s"&�>  uP� &9 u&9 u&9$ tX��SQRVWU����&�  �F �u!� E�N&�  �H��
 �pt�R�� �et�� �~�~ }sH�ʴ�� r@W��� &�}�QuOB�a�� �
_&�}�Yu&�E���F&�EW�g�� � [����~�Դ� rB�vW��� �y�� �� _���^S�� ���� �� _^�F&�D&�E &�D&�E�F�޴�i r,��	V���� � ^uW��� ����	 �q _� ����	 �d �~ hv'���. rW��� ���� �F _�^�_ �Ŵ� �J ��]_^ZY[XËN�7�W�J uW�w�W�A ^u��+�r;Gw����W�^� �
 [�� �~�Q�~��Y�~ð骋�+�- �ÿ Q+�AVWQ���Y_^tG��Y�&�6* �
��� u� u
&�<.uN� ����0N&8d� ���+؎�� W� ���G��_X+��������t�ڃ��+�s����+�3Ҏڇ���u۬�N���F��$�<�u���<�ul󤒨t����Ì�+؎�� � ���G����+�� �������t	��+Ўڃ��������t	��+Ў���Ì�H�؎�� � ���G����H��� �������t
��+Ўځ���������t
��+Ў����Ì�H�؎�� � ���G����H��� �������t	��+Ўڃ��������t	��+Ў���N���F��$�<�u����<�uk�¨� 6��S�Á��v[�PQVW��s�� ����6�>� &�=RBt� ��l� u$�h�6�>� ��(�D �� �N�� r���f �� �v � uD����2 �D �� ��x� s����D �� �G�u rW��� 󤸐H���� 󤫃��K ��8�t �: u0��2 �B �� ��N�: r��� �H���� 󤪃��K �_^YX[þ2��  �t	&�}�Vu��W�u6�>� �ˋ�3�&����_;�u����      @  � ���� ����PSQRVW�
 �v��
 �uJ&�  =\rA=w<��u7&� �� &�  ���� ���t���� ���u������Ы�ʃ����_^ZY[XÉ&H�L�J �� � �>CSu-�>sDPu%�>F�u�>$ �u����u� �u6�� 
��p  �����������RVW�øi� %�����Ȏ�.�I�&� 3��j�_^Z�>@�B.��=.�v�.�z�.�~��F�&����؎м 	�!��!��a !��B<��s�!��b�ȣ�
�J �6H ��V� �������� �������^3��ظH��� �ȣ� �7V�� � ��ȫ2���ë�ƫ�ث3����H��@������
� �� �^�L6�62 6�4 �4���Dt�6�6. 6�0 �j6�.& 6�( �4���t{���D �u�6�g2�L
6�F 2�6 F V6�l�7CC&�V &�vSQR��&�F6;6 v6�6 ��! &�F&�F&�F�ZY[��^&�v&�^V���؃�!�^�~���!�F���F����!���1���л �F��R��
����
�����:��
Z3��؎��� 6��
�E�� �  W��� ��@�	 �������� �������� ������� �D6��
�� �� ��� �@�� �@�� �@��  �� �� �B�� lC�� ġRB�03���3��� �F�d�� 3������ ��, �(&�D&�D&�: �m &�68 Z�.&�$ ���  Z�   6�F+�H� �� � ��(B�ں�������=�H�-�=6�&�6���6�Z6�[ 6�\ 6�]  SP�Z�w�X[�P� C�/<�uSR�C�/.��=�c�e�Z[X��X� .��=�� =  uM.�>�� u���r ����b�	 �����= �r-��r(�r��R��a �� <u�������- .���˜S3�3�P��X% �= �t� �P��X% �tCC��[��3Ɏ��� &� � ����������� �������� �������� �����&�� �SP���� ��
� �����t&;u���*�\O�\T�\Y�\^��� �\c�0�>�
�t	��
;Lu�DX[�3���&�  ��� ��� ����������� �������� �������� �����&�� �&�� �&�� �&�� �&�� �&�� �&�� �&�� �Ê�������PV�B����� .�<�����^X�                          ����B  ����        �           �                     ���NUL                                            ��         �� �D  �D  �D  �D  �D  �D  �D  �D  �D  �D  �D  �D  �D  �D  �D  ����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               /                    �  �         �                                  �    ��                                                                       �              �   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                       �                                            ��                                                                                             d                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               �� � ��EA�A��EEEIII�����O�OUUY�������AIOU��������������������������������������������������������������������������������������������� ��EA�A��EEEIII�����O�OUUY�������AIOU��������������������������������������������������������������������������������������������  �   ."/\[]:|<>+=;,                          	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`ABCDEFGHIJKLMNOPQRSTUVWXYZ{|}~CUEAAAACEEEIIIAAEAAOOOUUYOU$$$$$AIOUNN��?����!""�������������������������������������������������S������������������������������                  <�s�,�S��
�[�           Ȧȥȥȥ&   *   �P  �P                                                  l                                                             ����   �         NO NAME     &�O �              ��	
		P 
!
T�VR2	UW	S$&'Z�������� 
!
"2	#$��"                                                                                                                                                                                                                                                                                                                    �  "    2    �      �  " �    �         ��!>�  c:\wina20.386     6� �u6�6X�(�>  u7��
    �W�  �@  �@  �B  lC  ġ  �D  �@  �@      ��� .�.b��� .�.f��� .�.j��� .�.n�� .�.r�� .�.v�� .�.z�� .�.~�            .��.���#�y .�.�.��.���$�e .�.��(�[ ��? �.�! �Ћ��V�ڋ���' �!���&���F ��������X[YZ^_]�SP�.�cX[�    �   � ���QVW.�6g.�>k� ��t_^Y��SP��.��.�&��Ȏм��.�c�t.����.�&�X[�˴�<t2���2������<$t	�� ������p      "    2    �      �" p        Q� ��Y�                   \COUNTRY.SYS                                                    � �
  /  �  �  �  &  �  $    , . - :   �  ,           
A20 Hardware Error
$6�66�t萐6�66�t�QW�)��_YQ�<t�.�~.�|�ˎ���3�P6��&;E/X��3�����6�66��״�6�>	�� �t�G��
�t<t��_6�>6�_���<$t�������  ː����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      �mf�  �  �  �                                   �d .�.��Y .�.��N .�.��C .�.�9 .�.�/ .�.�% .�.� .�. � .�.$� .�.(�.�>4 t� s� ���5  SP�.�0�X[u����SP�.�0�tX[���P�
�uX��� �) &� � X��2��A�X�!2��B�X�!�P�k r��� u�D &�  <Zt��& @����X�P&�> u"&� =HIu&�
 =DDu&� =ENu&� =  X�&�   �  &� &�
 &� &� �V�R�!&�� =��t���^øX�!
�u�X� �!��!��
�������cox    �A  �         ���                 �    5                                                                                          ,                 ��  ��                                                                                                               ��!��!��!��!PSQ�ێË��J�!�>su3�> t,� �H�!r#��3�3���! ��������I�!�Y[]�H�!re��, ����3������>L! t�ŴI�!�b��&�  �������H�!;�r+�H�!r%P�+£`��X�N�O������I�!�� �����                                                                                    �9  �   \   l   �    /\�  j                                                                                                                                                                                                                                                                                         ARIFYNAbort, Retry, Ignore, Fail?reading writing  %1 drive %2
 %1 device %2
&Please insert volume %1 serial %2-%3
%File allocation table bad, drive %1
Invalid COMMAND.COM
!Insert disk with %1 in drive %2
!Press any key to continue . . .

Terminate batch job (Y/N)?Cannot execute %1
Error in EXE file
"Program too big to fit in memory

No free file handlesBad Command or file name
Access denied 
Memory allocation error&
Cannot load COMMAND, system halted
!
Cannot start COMMAND, exiting
.
Top level process aborted, cannot continue

� ; �     �  Write protect errorInvalid unit	Not readyInvalid device request
Data error!Invalid device request parameters
Seek errorInvalid media typeSector not foundPrinter out of paper errorWrite fault errorRead fault errorGeneral failureSharing violationLock violationInvalid disk changeFCB unavailableSystem resource exhaustedCode page mismatchOut of inputInsufficient disk space������		!	2	M	_	p	�	�	�	�	�	�	�	�	Too many parametersRequired parameter missingInvalid switchInvalid keyword $Parameter value not in allowed rangeParameter value not allowedParameter value not allowedParameter format not correctInvalid parameterInvalid parameter combinationA
U
p

�
�
�
�
�
Invalid functionFile not foundPath not foundToo many open filesAccess denied Invalid handleMemory control blocks destroyedInsufficient memoryInvalid memory block addressInvalid EnvironmentInvalid formatInvalid function parameterInvalid dataInvalid drive specification#Attempt to remove current directoryNot same deviceNo more filesFile existsCannot make directory entryFail on INT 24Too many redirectionsDuplicate redirectionInvalid passwordInvalid parameterNetwork data fault!Function not supported by network'Required system component not installedQbq������&A  Nj��������		!	2	M	_	p	�	�	�	�	�	�	�	�	                                                                                �  ���� 2Eg             ��<t��<t�s<t��<t�_����m�	rմM�!�k�y��t��t�4���t��r��w����� ���X�v�uP��!X���tR�uN��s@�nS��  &� �� t�ôI�!&� &� �I�!��u�[�n�� ���k3���{�|� 9vt�v���&��8ju�E��P3���
�t�.nXú���>s t�>v u	��o����,�f�>s u�� ��
 �� � L�!�v  �/�I�!��P�!�k�>j u3��j�.	X�	����ؿ� �@ �Q�!&��P���!�v� �j���>j u� ����H�!�
   ;�s�;�������ôH�!r��j �/% � r�/�;�v+Ё� s�/�!�/؉f��+�;`t#���w3�������N����Î`���`�؎м
� 3����x=��t�.�!�>v�u����;ht��&�r;ht�a��� ����`��3+��f� �.^��� �PS�ظD�!s��% ��[X���� ��63ۋp� :�t�>�!� C:�t�>�!�. ��� �>�!C���>��u�����/�� �SP�Q�!���4 �&�&� ���X[�� ��SP�Q�!����4 �X[ú����e�M�u���u���(�>  u	��!A� ������ �	� ø�!� �!�E�� =�!s= u���^�����غ�&3ɸ B�!r����`� �?�!�P�>�!X�r;�t����q���`� �S����3ҭЃ� ��ú~�"%�
 � �!�J���!�U���!������B�e��!��:It:Hu����
�VQWQP�݋D&�&���� ��
��XY_��R�Z�&mA���Āt
���u���j��t�s�>3UVRQS�Y�![YZ^]�>�2����s� � ��t��u��>��vB��� �/<�u*S�߸�/[r��׹��2����E�$�	�!�E� �� �>3�>������> t�]�1F���t���6����I��|�6����:�> t�������>uQ�6W��� ��_Y������J��mt�P�� �m t�X�� �mt�a�� �h�� �z�t�� ��!� �Y� �m t:Ft)���mt:Et��:Dt���mt:Gt�Y��e��t�>s t�N�p ���� ��L�!�c�t�d����
�t�>v t�v���> t�>u�| �>v t�v���ċ����Y^�
Ϻ���� ���}VPSQR�ދ�3Ɋ��� ZY[X^�R�ڃ��㋟
�����Zì<%u���1��	s� FI��д�!���SQ���؊�_��t'��t+�� ��������P$0<9v�д�!X������!��
�t��!C��Y[�P��/DD�=.t*= UtPPUP��F�F���F���FX]�X�3����uS��2���Ŀ�[�PSQRV� ��;t�Z ;�rZH���;>�rG�� �  � l�!r?�؋�3��� 3ɸ B�!r�5�@ �?�!r�u
F�5�u����>�!����&�=�u�^ZY[Xˊ�ȸ X�!���ɀက�
ٸX�!����2��X�!�      �
�P���!� 0�!=t�S"�[���&9 t�� ��&����£�!��
� ��/< t���/=��u���/��3۸��/�A
�>��
� U�/�u&�6�&&��&�&��&�e�������� ���!� c�!���6���� ��
 �� ��y������/% � s�/�!� �'�+����fP��&�Õ������J�!X��!Z ��! �������!+£`�, ��t�>�& t�����!���e�\ 
�t6�:�e@��>L! t �>o!&�}:t��� ��� �� �&�E���!�.!�k��� ���2���3ɉO"��!�O"3҉6Q"��!�O"=��u�}=  tHVP= u5���6Q";�t+�:�!t�<	t�:#u��b:�!uZZ�� :�!uZZ� X^�����z�떁>H"�!tG�>H"�!tT�>H"�!tv�>H""u� �>H"7"t|�>H"�!u� �>H"C"u� �>H""t� � �>z�u� �\��z��2��>s t� �G��s�~��>?!�u�?! ���>�! t� ����!�?!����t  ��s �6v�?!�p�>�! t� �����!�J"�������!���>�!u� �����!���1���,V�6J"�ָ=�!r`�ظ D�!�u�>�!�N2����D�!r��&�>�&t*Q� 3۴>�!C���ڴE�!�E�!�E�!�>�!Y^&��&�1�^� �n���#�&�>�&t�&��&�S��V3ɬA< u�6��!N�Q� �6�>o!� ���t�����+�6�>o!�� �O�q!� �>o!Y^�I6:�!t����Q�!� &�E�:$uFI�o!� =�!r�ش>�!Y^����"�?=A u�#�Y��!�>o!� ��َ�>s t.�P�ێ��!�
 �~��ث�J��ث�U��ث� �?�.%�!� �� � �p�����6o!�>L! ����u�q!W�I��_s	�q!�� &�>��|:u&����
�u�&�>\&�\&�&e��@&�& ��1��&�� �S����3ҭЃ� ���h�>?! u� �H�!r����!��!  ��3�����6��!��������6��!K3��o�!��t	+�sB����t�k"����!���;�!w��! �裍!�> u�� ��n� ��3�� ���3�����������
 �>! u��!�!�!�.!�!� 󥤺!� =�!r	�ش>�!� P�� �J!X�H!=A t6��!� 8�!r#��Ru-�  �.!� 󥤺.!� =�!r�ش>�!�M�H!=A u���J���I�!�  �n�  �<5�@!��&������B!�@!�>v u��"�������/�>�&t-�&��&&�6�&� ������&�}� �r&�4�����3ɬA
�u�á`�>btS�˸�&���������[�R��K�㋟;����Z�� r-�@��( �3�QVW��< G&:E�u��_^YtQ�" Y&�= u�����W� �W� Y+���à�!�2�� ��<�r,�S�����[�:�!r:�!w, Ã�V���D ^�SPRW�Ȏ؎��>s t<�/5�!�����>�& t������@�ظ/%�!���>�!u�C�>���>�!u� ��_ZX[þ� ��!3�3���!=��t2=  t���>H"+"t�>H""t�>H"7"t�־�&��t���g���� ��Ȏ؋���Cu�����3��>�&uSQ�3�!Y��r3���[u�ȃ�����������[����Ȏظ3�!��u�>��C;�t6�>�����J�/����4u)�4 ���ȃ����������뽱�������P��W�_�o�VW��>L! t�N+��� �>�& t~�tv��� +��tO� �M!�t� ����M! +��tO� �c!�t� ����c! +��t#O� �q!�t� ���>o!+�� �I�t���O��� � �>  u�L!�˃���������H�!s� ���tQ�+���+��Y+�W+��_�M!8tP� �8L!tE��!A�S!�\!� �\�u�G�!�	 �S!��;�!s� �\!��;�!r���;�!O�W+��@ �_8L!t�c!8t� �9o!u�� �o!�q!� ����L!_^��  ���Ë׿��&� �«�ë��ÿ� ����������� C�/<�u�C�/�0�2�               /DEV/CON       \COMMAND.COM   :\AUTOEXEC.BAT  :\KAUTOEXE.BAT �    �W  c3   PATH= C:\MSDOS C:\DOS PROMPT=$P$G   COMSPEC=\COMMAND.COM =az CKA            �W          �!  �!�!	�!�!�!�!"""".":"  F"N"    F"N"/P    F"N"/F    F"N"/D  �  F"�!/E �    �       F"N"/C    F"N"/MSG    F"N"/?    F"N"/K    F"N"/Y              Incorrect DOS version
Out of environment space
^

Microsoft(R) MS-DOS(R) Version 6.22
             (C)Copyright Microsoft Corp 1981-1994.
(Specified COMMAND search directory bad
7Specified COMMAND search directory bad, access denied
8Starts a new copy of the MS-DOS Command Interpreter.

8COMMAND [[drive:]path] [device] [/E:nnnnn] [/P [/MSG]]
*        [/Y [/C command | /K command]]

H  [drive:]path    Specifies the directory containing COMMAND.COM file.
M  device          Specifies the device to use for command input and output.
E  /E:nnnnn        Sets the initial environment size to nnnnn bytes.
M  /P              Makes the new Command Interpreter permanent (can't exit).
F  /MSG            Stores all error messages in memory (requires /P).
J  /Y              Steps through the batch program specified by /C or /K.
?  /C command      Executes the specified command and returns.
K  /K command      Executes the specified command and continues running.

LThe /P and /MSG switches may be used only when COMMAND is started by using
+the SHELL command in the CONFIG.SYS file.
F##�#�#,$z$�$%U%�%�%,&y&  8w5 E) �"�{��                                                                                                                                                                                                                                                                         ��!.������x=��t�.�!.��3�>v�u�&�����м$�������W��� ��6�᠀6�d���t	6����>r t�r �硴;�!�>� t
�>� u�(2�j �Ȏ�P�$�� 8�!X+�S� ��[�t���= v% ��&����nt��1r���u�|�u���u�*�>v u���u�&1��� �� ��!6�����t�u2�nt�t1r�|�u���u�!�|�t�6��� �� �� �{ ���tB���  �d��/<�t%���� ���u���� t
���  �]�>v t�6t�6v�f�3ɬ�A<u�I�e��9�	]�!�]��!�ᠸH�/�t�
�!��2���ᠿd���t)3���m)� �����d��L2���(s���,t��0�� �$4s�H��T����קu�>�� t߃>ڧ tؾf�����)�!�է�:u���߀�A<�t�>ا�= u����*��%�� �	 G�*������ V�f���(F���(t
<t:	�u�N3ɬ�<��O���ш� ^�>ܧ�>��6��u���\ �)�!���>秉>��6��u���l �)�!���>�> ��>ܧ��#>���>"�����%�
�u���9*�8+�����t���>v�t������;�<t6�<
t1��&�1�t#&�>�t�@t&���t&�&� ���Ëֻ �@�!�j��JS�;���8T�YNr���!��u��!<?u�&�1@�<u&�&1��$�:�u��:�uϜ�д�!���'��VWQPS� ���&�>���t�[XY_^ø ���3�&�=U�t
� = �r���&�]2�������〿 &�G2��u��؋�F�t�����<?t�< u�.�<�.�>:��뛻���H�!�H�!SP�"%.���{�!�ڎ�Z�U�!�ں� ��!&��, [��Ӊ ��J��B� �ځ� r3۱��ڎҋ�3�P��.�6<�.�6:�����`rÃ�t
��t�5 �.��t�e�y0�{�B�����Q���E���Q�����Q�. ���  �-�>���%��#��%��%�>��'��R�c�!R�c��!��!� �!�cZ�!Z��o�d�u �c��>  t��&�f���%��A��f��؎�6 �6
 ���\<:YZt1���t8<@u�o �-�� �
 � B�!&�M���3�������u���wA�f#t��sQ��hA�
��� sD<%tJ�<u܁�g���&�e��I� �>o t�nut��>�t�:%��f��%�,%�<t� ���<%t�<t�,0r9<	w5������&�w���u�m��I�<tA��� s���2���O�IW���0���<u&�E� ���_�r��I�<%u�=&�E����Q��!Y��_r�o�����u��t<u����&�/�I�!�������H�!S�H�![&�/����%�u��% �u#��% � r&�/�;�r��;�r+؁� s&�/&�!���،�+�S� ��[�t���= v% ��&�Î�&�>�t�)�h�&�>�t���-&�n$P3�&���t&�&�>�t��&� P&�>�t�&&�� �-����/�N�ֹ �!�Z*�فÿ Q���S�H�![r$P�  �˺�������;�r;�wX��� I�!� X&����ZX&�&�&�   &� ��3��|&� ���t�}�| &� 3��}�n&� &�  &� &�
 H� �߹
 ���f��
 ��"<t�&�?�����"t�<t
�����I��2���]���J�!�>v�u�v��X�n�;�ZXX�#��#��%��%� �&PS.��.����tB���nu�o &� �n&� �}&� �|&� �I�!��&�3��[X�P�A��� r���
�u�IOX�SQ�d�t�� ���u�� �&�>  t� &� &�
  �Ȏ؋M����u@�O��Ȝ�y��?�!s!������S��M�f��g� ���j��� �o�3ۉM���O�C;o�r����M�<uu��&�&�>  u&� �o���N�
t&� ��&�. t&�> t��5�
�0������d��d t�f�3���>v�u�> u�v��Y[�X����$���>� t�7(�� �!�  �� �� <tՋ��� ���G�7�u�&�%G:�t�� :�����GG�u۬<t�� u�� �����!��V3ɬ<t�� tA��<=t<t(����<=u �x <t_�tN�<t��<t��i u����:�L���\ u�2��-��R u��>�� �!� !��է�4,�� � N�!r2�������t��
�t��� �΁� (� �� �e��f�������{��k��|��
2۬<t���t,0����Æ������&k2�:�s���듎���uÎ��ؿ �u�	 �=�t�5����<u��< tۉ5����t
�Y��{t�����VWPQ�f��c���f��| �YX_^�������>� t�|&Î����t�3��� �
 �  �c��] � � �uA����&�>��z�r<:t&���<
u	�j�r<:t���u��w �� ����V"�K�r�] &�>��Q��Y�t&:u�GI��Q��Y&:� &:u�, &:u�G���p�&�>>�}< w�<t�]�<u��V��&�  � �.�y���r�>�!�c ���  � =�!r� �
 &�y��ظ B�!&�M���Ë����Њ,@�����t6��&� �� t�ôI�!&� &� �I�!��uԈn�  ��&���>v �u�> u�v����nt���t��3��ơ}�؎���� �!�>E t�G�G;Iڸ  �r)�O��Gu�7�(8D�uA�:8Du��+ʃ>E t�Gu�O�Q3ɸ N�!Y�� O�!���r�  �E�u��7�K�>E u���< t�u�2��3���3ۿf��D�6K�  ��(�w	F�F<%u84uFV�K��
���OA^��I<u���&�e�&���nt/�>�t��� W�
_&�E� �%�f�����G&�E����� ����H�+�e���&�>| u�&�>� t�#3��� r�<%uۋ�
�u��� r�%��=INuǬ
�u��� r�<(u��� t��)u�J���OF�� r�=) u�5������w���)8t� r����� =) tG� r�%��=DOuЬ
�u��t r�PSQRWVU�:�� ���*�&�}�9��]^_ZY[Xr<&�6}IO&�G&�>I&�D&�E����&�&K&�|&�>v�u&�v ���#��%��%� ��B;��}�ڸէ�P'�7�����������>v �u�v���P.��&�}�t���I�!&�}  &�| X���
�� �� �s� �C���� u
�3�./�����>���!�\ G�?� ��rE�>� u>����� t
��
s�&����?
��rI��� t��r<��� uR�7��t��F�� u�� t�`��#��� �#��%��%��� �>%�u�%� ��� t������ t�ÿ���>���*������ 3�������C�������������r�U=��t�SE�#���g��AEþ� �;=��t���ú$�� 8�!r��t�e���� �ӿD��!s�D� ���� t�&������ t�&����@ �ؠ� 
�u�2�������D� ������!����/��.���� t�.��>��:u
���$�,@�\ ��#u���V�6����������� ^rtA�6@��/����u3�>>� t���%�|:u��<..u�| u����\ �)�!�����#5�!�I��K���#%�!���� �� �+r8����s= t��8S��[��� 2��S�����[��  P�..P����XX�r���]= t= t���S�t%�>\�.t�\����v�\����s
�\���� �þC�3��
�tFV������.��Nr������Ї�^t��Zi������������ ������	��	� �>D�u'US�E��/CC3�&�G;�s׋�&�;�s�;���[]��&�Ë������� ��&��Ë������� ��&���&�G&�f%:��&�G&:F������� ����� t3�e���d���B����� t�C��A��M��I����7��;��3�����6�\ �!=��t����.��0��s��B�Ë����>��2ۆ3ɴN�!�r�S�@t3��O�:���II�x����ø`��w���@ t� ���r��3����r����Î�3���p r���v r�]�s��� ����&��Ã��� P��* P�*.P��P�Թ �N�!r,���� �O�!r������;= u�~ �t������
�t��������&�<t<�t�Ã��������Lr��� ��
����� ���U ��[ �U ��!��r��U ��!��r�Q��&��"�"&��:�u��3��1��3��5��A��I��K��>C� t�6 s������r�)�����r����= t= t���>1� t�I����3��&����i�r!�  �x�r�&�+�= r� ��&�����@�þF�2��� 󤬪��
���ȭ��u����� u3�����t�̱��
Ī�3����Ȫ��C� �Ë����� ���� t	�����!����V��� �w� �
�t1<-uJ����� �u�у�������� ������������^ÿ��3��a=��t=  u�ڀ?t� r���� ���VS�w�C��
�u�C�C�C�;2Ҭ
�t4<-u������� �u�ك���u���
ʈC����s��[���� [�^���V�w�
�t
<Ht�~������^�QW�G���� ����.���_Y�dLdddddddddd]����>��$���
�u��>��;�!�W��2�������_��V�w�^����1��7�u�9�&�G&�W3�5�;�=�Ìَ��.��tD��� t3��>����  t���
2������O&�}�\t�\ ��%�>����>� ���.���؎������ � ��A�ы����6���  t���
������ � ��t!A�B�.�
���	��.���  t�x�
������� t�<��$� ��� t���B � ��� t�"������� u'��� t�c���� �?
�
�l���=���J���������o�� �� �� �2�����  t�o����%�o����=Ã>1� t�>-� ~����m=�����.��-��-������&�Ft����F=��@t���9=�&�V�!�&�V�#��ޘ�!=&�F�tH��% �Ћñ��$������2��P��dr��d��?��A�&�N������������J��:���<�����&�G<�t������$�&,��-�����<���� uG�'� �1���� t$P�A��t�K��I���&,��-��Ù�n<� X�*��e��a<�V��[<�{ ����Gt�[�����Gt�]�� +��� ������� tSQ�:���p��<Y[���H�/�à\ 
�u����@�:ø	 �#��%��w�6%��'��%���/��>/�w��ÿ7�� 2���PSR���Z[X.�.I�<Ar<Zw �W����
�t������_��@ �؃>J (u(�&蘿��

�&o���&`���a�

�&}���~��&��@���o�@�`�@�a��}�@�~�  ø���Q�����\ 
�t���� ���J� �/�u��Àt��SR�J�ӻ �/ZY�ut����:�t�ٿS���A�:���I��
 ��2����ǳ
� 2����0�ઊ�����S��ERV� =�S��!s�EBL� =�S��!r�Q��ش?�@ �c��!r;�t�m ��i�>�� t��S���@�!<�u�p�����&��(�= �s���  �������������'� ���������+�% ��&��������������ËQ����t�>�!�Q����(��&��SQR���3ۉ?��E��G�= rz=��sM�Jrp�,rk��sg����� ��CE��G� �Њű��% K;�s�Ê��2����2�?���� r*멡?�A�C��G��E�I�K�M�O��	 �3�ZY[�VW������2�����8 P���t#��3ҋ˻
 ����ыϋ������ыϋ�� [��<
r��2�_^��"VW3���+��r���� ���ыϋޓ��_^����3ҋ��+��r�؀>�� u����&���������&�u%���ٱ���=�r݀���؋�+��r������&�&�_�Ë�+��r+��s��PQR3ɀ>�� u	��������$��������Ëء��q��&n��ы�������8 r1���@�&n����3�������������ы��������� s�ZYX�SQ�ʋи B�Q��!r�?YZ�!r;�t�ú����7�2��aþ� ��  �~�3�3��=��t>=  uh�>w��tV�6y��|:u�| u� �?�(^�̓>� t� ���5����s���=  u�>>� u�>� t�	�� �#��%��%��l�� � �3�3��=  u.V�6y���^3��=  uV�6y��:8Du�#��%��%�
 ^�h�l �)�!��6�^� ��<u��.�6�t�s���=  u��>>� t�|��6��T���t,��\ �!<�u�5P��P��	X��t�X= t= t�K��3��þ� �l�3�3���=  uV�6y��^�l���t��9�B�t�T��� l�  3ɺ����!s��%����'��c�ظ D�!�t�s�����B3ҋ��!�q��s�� B3��!�#� ��3�.�>#� t�.�&�.�>s��t1.�>s� t.)q�.�s� �.;q�v.�q��c.�q�  �.)q��?�!s�g����H3�P��X�=  u�}�u
+�I&�#�S� �@�![r;�u�z�I;�uû � D�!�u��
þ� �Z�3�3��=��tE=  u
�Z�3��t6�lW� ��/
�t#���/=��u���/�������3۸��/_�����	� ��U ���3������G� �?�>���!�U ��!P�\ @<@u��A�8�X
�t� ���o��׾F�� �2���.�R� i�\ ����!Zr�4� ��G��4� �#��%��%���SQRVWU�Y3��!]_^ZY[þ� ��3����=  t
��=��t�xS���? ��[
�t4�3�!��<v��A�6��~��04���r	��r
������������4��0�!P2�2�X��2�4�����3�r&�= u
�i �>�U �8&�G
�t0<$t�D ��&�G��
�t���X:t�? u���W�W_��ú��3�=���
�>��<��|WR�д�!Z_ô�!A����2Ҿ>�����A�:��
�����>%��G�!��s����N3�� �>��%����=3Ê\ ��@<@u���P�A��G�!s�	�>���X�:��
���2��3��O�Dt`<;uF��<t4�`t������<;t��u�<t< t�<	t�%��%� �#���
2���q�E����3��< t�b��3����T� �#�&�= u
�z��2��������� t����� +ч���a2�� �/<�t/�D� ������!r����𡚧���>� � D�!�t��u�R �,��<v
<t� ���@ �؋J �6� 
�u���� �����R�3��Z3��ȴ�2�����3��þ隬��2�����!����� ��3�3��1=��t=  uV�6y������< u�^����t�����=�!r�ظ D�!�u�>�!����o1�@R����S�R2�ָ @� �![Zr�2����D�!S� 3۴>�!C��[�E�!�E�!�E�!�>�!��� �p�tP��� ��3�3��i=��tc=  u[Q�y�����Y���7uH�� �/<�t����9����f��!s@= u�Y3��!= u���������Y3��!=A u����������f��!�������0��� �u�3�3��� �3�=��t=  u6�>u�t	�� �.��)V�y��@��:.�� �^�V�6y���< u�^�u�� t�_�3��d��`�!s���%�3��'��B�%�d�����0����>s t
�>v�t�+ٸ.��>����/���&�&� &�&�
 &�&� ���I�!�L&�k�!3҉6���/<�t	=  u@� É6���/<�t=  t� ��#��%�� �%�= t�6���6%��'�F��� �V�^u��}�V�S� �t�3�V�<t<=u��À<u�����^��t����MS� [��t��n���<V���ǜ �虹 �u�ǜ��^V�<t���^�>ǜ t�������3�&�eP��GXu�|:u��c,A����&�e@&�>�&� ����Ot<t���2���ǜ O&�>\Î��3��< t������
�u���g.��ܙ���V�, r���� ��&�< uN�p+��^þܙ���� r�� ��A ��&�3�QVW�� tN�GG&;E�uI���� G&:E�u��_^Yt�Q�d Y&�= u�����W�O �W�M Y+���À<t���F t	� �� ���b � <=u�þ� �
�t��O<Î�&�3�&�= t�� ���=�2�� ��VP.���6��< tXP:rF:vF��3��3�@X^�<�r,�S�������[�
<ar<zw, �QS����R �ك�;�r?PQS�2�[���� �r�����C��˃� ��;�s�J�!������YXs�<���&�  [Y�P��H��&� �����X����>r t�硴;�!2��þ� �u�3�3���=��t=  uP�>u�u�u�3����u?�=���V�6y��^�u�3���u%�3�B�u�;�!s����= t
= t� ��`��C,��? r9�9�!s���= t(= t� �!�3���!�N� �!r�H���t�S���c��,þ� �l�3�3��V�=  u�3�WV�6y���< u�^�l��$�ZtԺ%�3������ru�:�!s��:�= t
= t�	 ��f��+��#��%��'��%��%�ÿ硊�@<@u�����&
��:����G�!r��R���k+Zì� t�N�< t�<=t�<,t�<;t�<	t�<
ù �< t����< t��.��Ī��< t���2��æu��|� t���P�QW�������E� �%�����*�E�r_YX����9�&�>� t�]	�����P�/8&	�t</t<\X����  �\ ��r3�v�B�u,�;�!s��= t= t���� �]�?�] � �2��� �6��N�D��>ԧ u��td�΋�R;�t����tF����u��J���Z;�tV�΋�;�t�ԧ ���t�F�ԧ��P�.8Du	8Dt�| Xt�D�<:t!�>ԧ u�4�u��� �;�!s �n������Ê���u�2ۆ\�;�!r�\�F�6@���>���t�\ �)�!�Ó�3��T�:	�u�� �F�F�<t�F�>����� �u	� ������Һ����
�t��3t)���� ����������������W���/�>�� u� �2�3ɾ���G�:��u��������G�GG�GG�u؀>�� u�z��"�%  t&��t�>��u��  P��t	P����(X��X����t��
�<�u�G��j��u�/ u�#��%��%� �� �����>��� t�����W�� �� ���2�.�	�< �_��5t���.�� .�%�.���.�9� R����`�Zs.�9�� �-�� .�>9� u���t= }����R����I�!��&�j&�r �-��5�P ��\ ���R �5�� K.�9��t�jՌ��Ѽ
.�.��H���'�	�3Ɏ��f����<"u����<u�Q����*�t��=  u��D�  ��<"u��t�<"u�����<u�Y������t�G��G������<"u��t�G���<"u���<>uW8u�&�����<<t<u�&��	 � W����Q�M �<t���t:	�t<"t<<t<>uN� Y�a�����Y�T<<u#����<>t<u����	 �aW�����뫊���|t��|u=&�>� u&�&n&���a�<t<|t<|u���:+߃��t&8E�uO2��_�%G��t����&�>� t��&�>��f�����<u��e�&�>� þf����6���� 3ɬ�<tA���� ûd�������� ��/< á���6���B� �>� �6��������MQV�Z����[+�Yˋ��ԧ �6I��r�tIF�ԧ���!�u�>�<?u�B�<*u�B��|�t:	�u�N2��F<u��6�����þ� �
�t�� <ì�M�u<;u�N�RPSQ.���>� u�{�u�	 �N Y[XZ�.�>�� t����� =���!r�ذ��G� �� =A t��=t�?��h�.�#��%�.�%��X��>� u� �>� te���=P�![rP�ظ D�!�u_�B������!� ?� �6��!r+;�u�>6���u7�B������!�+.��� B3ɋ��!�= �u�e���3ɴ<P�![s�U��ذ��G� �P3���A
�u�+�X�s��SQVWUPR�Y�!Y[�K�=A t�Ë�]_^Y[������VWQ���3ɋ�W�< t�A�����_����>��Y_^�.���>v t�>v��ð���r�R.�����A�!�9�A�!Z��� ú���������^�PR��������#ZX�=A u����͎���WV�;���r�������� C�!r�� u�^_s�.�&��&92�&��&:��3ɴZ�!s냋ش>�!�9�Z�!s�q��ش>�!����6��>v�u�v ��-�&n��6��<|t<|t� �� =�!s�2��ذ��G� �f�3ɀ<u���|8t��<|t��u�t�AA��<t<A<|t<|u�&�E�I&�e�N�6��Q3ɸ <�!Yr��ذ��G� ���&�e�N�6��z�������>v �u�v�����.���Ȏ����s#�$�� 8�!��  �d���e�� �l ˾� �6�3�3��@"=��t=  uG� ���ӗ�՗�×�<"�� =��t)=  u%����6�����QR� 3���!<�ZYu	�+�!
�u�������"�þ� �H�3�3���!=��t=  uN�#�,�!������������!�� =��t-=  u)�.������6�����QR� 3��!<�ZYu	�-�!
�u��"����!뿎��&����P.��2���
�t�.nXô,�!���.�1�.�3��,��L!ø 8�\ �!��.�
�Hx.��t.���¶��".�6䗺ߗ�!.��  �
�d�� �x��!3��q����f��6�3�3��� �3ɺ���� �
�d�� �M��!3��F��]��f��H�3�3�� ���< t�<	t�Nù��2����W�_�ѿ�WQ�Y_���9��PSQRWV��)� �����3��D�է��������  ���  �f����>| u���2�e���󤾙���� �6��3���� ����:s	�t� ��)�� s�������^_ZY[X�SQRWV��f �>��@}O���������է� �G  �O�w�6��76{�+��w�6���w	���>������}+��� ��>����
� �� ��^_ZY[�PSQW���t�>���t����է� 	o	.�������������_Y[X�P�ó��[Ó�SQRVWU��קt�� �[���� �!����ʭ�>̭�>έ�� �-��r֋�������tk��-��6է�ا+δ:��r8dt��A������ �Ѐ�`�Э���r
�I:ЭtANV��� G�!��^�Э�= t	�= tG���8uFI��� �קu�;�ا+է��-�� ���u�s�3�� �-��έ�6̭�6ʭ&�|.u;&�|:u4Q&��&�D�E�Э�EV&��� ��`����� G�!���N��^��Y+��6ʭ�����tI��I��w��Э���O�Э:E�t��ҭ3ɬ�
�u��ŝ]_^ZY[�P�/��t�\�ЭXâЭX�SQRWV�������6έ�6̭�6ʭ2ɬ
�t:�t��t�����2ɪ���6έ��3����t!�Э
�u:E�t���
�u�����}�� 
�t�����^_ZY[�QRWV�R���߭3Ҁ}:u���߀�@� G�!ZrL� � N�!rI�ѭ �ҭ �E :ѭ~�ѭ����ҭ� ��<t
� � O�!sڠѭ�>��t����ѭ�
�����  �^_ZY�WV�  ���� ��u6������ǧu�u� �#������u�u� �������u�u� ��  �>��t=  t���� ^_�PSQRWV�����է�>ا�= t@��ڧ+�A�.���	��� � ��+ʃ�;�������>��u
O��?���� ������^_ZY[X�SQRWVU���S��� H�!rD�����D3��է���3��էI|$������է+�&���ا+�&�W��ާ+�&�W	����������]^_ZY[ù �] �<?u���� u/����� ���x �
�!�
�t��*��s�< t�<���uѴ�\ �!��t������R��Z�>%�u�%� �w�������!��\ �!��tӾ���ˤ�
�������>��ڀ u�G �%�����ˤ�%���������!�s�< t'<t뼴����!��u�X�= u�g��=�����a������!��\ �!��t�y��-�= t�V�����6��� r��u�nÀ&n����� t	�� �m�����n������"�b �3ru��!�2��!À� u�2��!�ں�����
�u���R�ڭ���*���7Z�2�  �� �.r
u�!����!À� u��T�!�غ��뽾� �< t�<	t�<=tN���3�3���=��t0=  t���'�>v��u�
 �3�
v�����3��=��u����ȝ�i���W� ��#��%����_ÿ���*�!�QR������Ρܗ��W�p_� � �ZYÊ�2��#e�!�3��'��W�����$��*�� ��{��@��%��?�����B�����Y��>�����硢Z�������b��d�����j��f��h��^�����������"����`��[��_��1��\����������w��x�� ��C��������>�����a�H����,�����>��(�� �+����)�3� ��6�����a��ǀt�`���u� �� t�"� t�� @��@ t�"�@ u�"�� t�� @�v� �ŀ t-�<yt
<Yt�� @�� F�"�@ u�"�� t�� @�v�	. �	."���#t
�� ���6�r5�[��r/�ǀu��V�{�� �+ƿC�ǣ@��?�A�>B�� �  ^�)��>`�u�>�u�>a�u�N����`�������Y���
�u�%��%� �<v�%��%� �#���>�<u ��A�:�F�C��� �  �F�F  �F
�~u�:8D�u�N�E��F  �*
�~�= u�`��:8E�u��F �N�
�"�� t�T�!��2�x�.�!3� �+� ��
��u�	. ��� u�>� t�_��>�D � �E�W��61��6'�������>� uC�#��%��%� �%����'������>� u3��$��*��%��6W��硽����6��À>`� u�3�6W��+� ��{	r��ǀt���u����>��u������� �\ � )�!�< u�����:t�@ ,`�\ ��w��V�t�P�2��,�
�t� ����>��2��Z��>���?���>v� tq�����3��`�!��u�>� u�И���]�N����>$� uB�Yr�>� u6�>w� uF�-�>�� u�>� t�%����� t��>x� t���%�����>� u���t	�И�o����� �>� u
��r�$� �>� t�2����t�� u^�%� �.��>���t�6W��6������3�6W��+� ��#�ǀt2��u��]��7迿�� )�!�������>���N�>� t�Z� ����Z��A3��$��*��%��6���6W�� t���������u
��P��>��!X�\ �!
�þ���3��`�!�� � l�@ 3ɺ�!s��؉��� W�!r
�b��d��(����%����'��Q�>�� t� �>$� t�b��b����� D�!� ��t�>[� t����I����&��*�+�u���>^� ue�&����?�!r����Q�>�� u�>_� t�ы>*�����u��A+ы�*��*�;&�r��>^� u돀>�� t�>� t�����>�!À>%� u�� ��t.�*��\t��3���� �*��Z� �\�*�r= t
�2uփ>\� u� ����d��b��>Y� t1�,�!������������
�Q�*�!����������������� 
֊�Y�� ~7�W�!r�B3ҋ��!М� D�!R�>�!Zs	��` �, ��u� u� ��1��%��Ë����� �1�  ��C��A�!�V�{�� �+ƿ��ǣ�����A�>��^�������À>�� u����%�C��'��b��w� � C�C��!s� �w��6k�� �DC��\�D�D�D �D	 �D
 �6k��O� � ��2��3۸�!< t�<t;�؊и e�!:�st:�st:�su؊�S��s�@� � ��s�!�@��s�![븀� t��׸ e�!R�.� 3ɶ�2��Z:�st:�st
�v� � �����v���&��6A�� �: r�! rG&�$�<Yu�v� Î�&�>� t���&�= t&�=/tG������3�2�&�= tQV�^Yt	Q� ��Y�����à�P� X:���^� �>$� t� �� u�>�� u�>� �N�u��Z�� l�C��! 3ɺ�>Z� u��!s�1��%�C��'��� ����$��ظ D�!����t3� �$u	�_�
[�tz!�t�D2��� ����!�� �_��Y��>Z� u$�>��t�\u�>�� u�Q��L�*�  �^�Ë��3ɇ*����\��>Z� u53����@�!�9�s�N�+�t�����t9��� u
�>Y� u�It�����#3҇ѸB�!�f��h��>� t��@�!r_�j�����%��>$� tH����� ~3�h��f����t!� B�!3ɴ@�!�>j� tA�j��@�!�>�!���>�!�C��A�!�$� ����$zP$�[�X$�_�Y��_�
�À>>��u�硽>��� ��2����
�u� �6@����� )�!�< t�?��S��C���:t�@�_� ,`����B��&��%
�t:�u�>`� t���2��4"���
`�������Y��>[� u%_�
�u
�t�*���3����uO�>*��?��>� t�������>@�� �<?u�< t�C��� 8t�.��<?u�< t�C��2����FuC�Ճ�W� l�@ 3ɋ��!_s���= t#= t= t��֋ظ D�!�>�!�uS�FtM�V�� t��:t�@�� ��`�z�s���֋Ճ��~����u�v�:8\�u�F ��F N� ��u�F  ���;�!r9��3���I&�G
�t2��)�t�G����O�
��F 
�u:E�t��F �N�t ���= t= u`�F  �~��t��F �v�< tK�.8tE�:8\�t�F N2ۆ�%�;�sVQ�΋���t	�;�r�Y^�;�r�Y^:\�t�;�!�s��������Չ~�F�?.� �Ī�ı�2��þC�����`�!�3��������3��>{��~������W3Ɉ����y�u< t�<	t��
�t��ǀt����-:�u�π��<u�:	�u��:8u�>)�u�)��\��X�>{��}� � �>{��}� �>)�u��uP��A�.�:�)X�>{��}� ��t���x�>)�u���<.u	�~��}��<?u��<*u0���>�� u�$�x��>~� t��?*&}�r���	���� ��������u!���>�� t��uH�>{��{��}���~� � ��g�t8<t4:	�t.:�t*<:t�_��>)�u�t ��F��M��6���`���N_���N�Q���� ���F���t�E ��A �� @�4<u	� ��� @���+ ���WQ���� �� @�u����� ���Y_� �_��êA�}��.�`�  .��.�&�.�6��.�S�.�U�  .�h�  .�Y�  .�%�[].�'�|<.�)�>+.�+�=;�	s���S&�&:s� [�#.�6b�SWU�j�.�a� uC��
r<�w	t7�	u.�a� u�?	�&.�a�AtN�.�<=u.�a�C�
sŬ.�C�N.�6W�.� .�f�&��6j�.�</t6.�<"t.�a�uT&�G2�.9S�s.�S���CC�&�� �i.�U� �`&�G2�@���&�2��tCS&��� [sACC��.�U� �4&�G2�@���&�2���@�&�2��tCS&��] [sCC��.�U� ]_[.�S�.�U�.�6W�.�Y�.�[���P&�� u.�S�.�< u� u	.�U� �P���� X��X���UQ&�O2��t�o	�s� ����.�.h��Y]�&�~  tE��E�.�a����rJ.�&a��P.�d�+�.b�X.�6d�.�< u&.�|�:u	.�U�	 �&�? t&� u.�U� �	� ����
P���� X��W&�.�>Y�&�&�eP.�h�&�EX<u
&�U&�M�Z<u&�U�P<t�<t�<u&�U�><u.�b�@&�E&�]�+&�u&�MP&�Gt��	&�Gt��X&�Gt�� _�.�.� P&��uPSRW.�U�	 ����[�_Z[X�0� t.�U�  �.�>U�	u� t.�U�  �.�>U�	u��o�� �t.�U�  �/.�>U�	uW� @t.�U�  �� .�>U�	u@� t.�U�  ��.�>U�	u&� t.�U�  �.�>U�	u�  t
.�U�  ��.�>.�u.�>U� u.�U�	 X�PV.�
�t<:u.�| u.� �	��sFF��^X�VR��.���r
�t� .��FF��Z^�<�s<arE<zwA$��=SW�> ���t�>�.8tPQR�e�»��� ����!ZYX.�].�ECC,�&�_[�P.�a��.�&a��.�<+t
<-u.�a�F� X�PQRV3�3�S.�
�tB�� r92�������� r,�ڋ������� r����� r��� rՃ� � rF�[� [.�a�t
���҃��� &�w&�< u����t�F&�< t`F.�a��u&;Lr6w&;Tr.&;Lw(r:&;Tw �2&;L|&;T|&;L
|&;T���	��u�.�U� �����&�$�.�U�	 ������^ZYXÜ.�a�u�Ýp����<0r<9w,0����PSRW&�&�
�u���L<u?G&��	��@�&����@�&�GG&�-�2 s����u�.�U� ���&�e��&��.�U�	 ����n�_Z[X�PURV�.���r<��.�a�t<=u&�~ uq�.�a�t<:u
&�~  u\F�\&:F u
�tRFE�&:F uEF.�E&:F u:FE�.�a�@t&�G  t&�~  t"&� t<:u	&�~  u�< u&�~ :t��.�6d��^Z]X�PQRVSV� ^.��  .��  .��  � r.��
�t� rn.��
�t� ra.��
�uY.���t".��
�uG��.��
�u=��.����u���.��.��
�u ��.��
�u���ds��l[^����)��[^�����.�U�	 ZYXÍ6�.�<�t�RP� 8���!XZ�QR3�.�
�t<.�>� t��u<:t0<.t,�<-t&</t"<.t���r� ��
 ���u�r�F뽊���F�����ZY�PQRVSV��.�D^u�.��  .��  .��  .��  .����o�r].��
�t_�b�rP.��
�tR��S�rA.��
�u6.�`�u;.�6W��|�,u0�D�..�`�  .�`�.��.�&�.�6������r_.��
�uW.��
�uO.�`�t<wCu2�.�a�t<tr/<w+��.��
�u!��.��
�u��.��
�u��[^������[^�����.�U�	 .�� ZYX�PV.�F
�u�.�D� <pt<at<mu$N.�D� <pt<at
�.�a��.�`�.�D� ^X�PWV.�>b�.�
�t�_ u$.�.�^.� _�?^.� _&� u2.�U� �)XV.�
�t�- t�hsGFGF��.�[�.� G.�>W�^_X� t	P������X�SQ�%��	 .:tC��AY[�PR.�
�t8�r,.�|:t&� t.�| u <ar<zw,`�д�����.�U�	 ZXì�" t�O u.�a� t�.�a�At	N����N���SQ<t)< t%&�}r3�&�]��&�9 t3�&�	C&:t��<Y[�SQ.�[� .�&a��< t6<	t2<,t1< u�< u� F:��&�}r3�&�M�t� C&:t��< Y[�.�[�.�a�u.�a� :���.j�;�t</u�P.�G����r����X���</u.�a�@��VS.�>^� u'PQRWU3��޸ c�!���]_ZYXt).�6\�.�^�.�6\�.�^��< t:r:Dw��FF���[^���������� �� ����1� ��1� PSQWVR���  ��P���2�X�� ta���WQQ�޹ ��Gt
�G  �G  Y��YP�>#��t����%�3���X_����Q� u	�Gu�O����Y�ށ%�u�%��W�1��$��6#��$� �#���Us���Z^_Y[X�>�� u��>1�u�l������&���t�ݺ����#��%��%��6�S� [�Q� Y�PSRW3Ɏ�3��.� �/�9��>7��.��/�A��>?��.��/�Q��>O��.��/�5��>3���=�1��>/��M��>K���=�E��>C��.��/�Y��>W��r�
���$�w�  �y�
 �<=�>[�� �r_Z[X���
��PV� c�!r�6k��m�^X�PWU� r����t���]_X�VS3�3ɀ��u��[����%��tļ?����= r=' wļK����ļ/��Ã��u���u���w����� 3����� t�T ���r�u럜��u)RUQWP� �/<�Xu	�ظ�/��s_Y���� ]Z�����[^�WP���2����IX_Ã�u�>W��t=��uP�w��W�X��W��3ɀ��t&�M�	.85u.�M���s-��t���t&;�.;u�	It�����r����u&}r2�&�G�q� �PSQUWR��o��6t�����t#�u�/ ��rZ�_
�t�%�����_Z�r]Y[�������PSR�o����u�, ��w s�Y�  �!2�������t;�t� ���rZ[X���u�&��!��� s&�U�!����t	&��!GIu���WPS���ٰ��u+�K��[X_�3��tO�@�׃�u(�!P&��Z Xs��@B�!�&�=u��������UQ����Y�!s�;�t;��u��]ø' � �À��t�ƀu�>r�� � ��W�>k��t&�= �t&:r&:Ew�GG��_Ïu�3ۓ��6y���6y���	v��7���0RA�u�t9��u�|
,u�6��A�"��u�|
,u�6��A���u�|
,u�6��A�3��3�3��6u��3��t!�%� &8%u
&8et:�u&��S�sGGBIu�V���t3M�>w� u+�D0&:Eu�<0u�t4��>t��uBBIIOO����W+��
�_Ys� Q�ʀ| t�tIIGG�^��u^�	���u3��tdUWQ3Ƀ>w� u;�Du�|�Z�(�Dt�Dt�Du�|�h��Du�%����R ��  rY_]^���
��>w� ur���w�  �3ҡw��y�
 ��X��{�C��@u�� ��u�
��{�CC�� �3ۀ| uǇ{� -CCƇ{� C� ]3�3҈q��D	:�v*����D�t�D
��{�C��@u�| ��u�| t8Ls*L�ъL�t$�Du�Dt&�G�X��{�C��@u�A ��u��D�u
�t�D
��{�C��@u�# ��u��Du�Dt�
�t�u���u�� U�QW��3ۍ>{��t�r_Y�����]�D0u&�PA�Z�s&�EP��&�
�tGA��+�U�]3�3��y� 3��D u$&��Du��tC$�y�
 �Du�y�
 �T�Du&&��Du�ĀtC���y�
 �Du�y�
 �(&�&�U�Du�ƀtC���y�
 �Du�y�
 �D@t)PR�82��{��!s���,�D
��ZX�D
,���ǈD
�����t3Ҳ-RU�]�y�
 �s 3�3��>{� u�} � �6��A3��D� �6��A�D�t �>{�u�X �g �6��A3��D�Z �6��A�D�O �>{�u�D�B �6��A�D�7 �6��A� �, Uô8� �{��!s�{�  ���-ËD�Du=c v�c Ï{��q����I:q�u�0 PAA�6{��]�y�
 �z �Dt�>�� u�D<|<~�aPA��pPA3�3��D t�D�e �6��A�D u�Dt�D�N �6��A�D�C �6��A�D�Dt�>�� u<|,< u��W�Uô8� �{��!s��� ���:���.Ï{��q��-�I:q�u�0 PAA�6{��QR���v��$�������!��
�t���s�Ȋ��!����� rZY�����PQW��3�&�&�&�&��&�C�� �� �!�_YX�PSQR�O �irA��3ҋ�B&�  &� �u&� ��&�  & ��&� ��&� ��& C��<Zu�� ZY[XøX�!��&�A�X� �!�3����A�X�!�W��� t�</tN��-�$�<Su� ��&���<Lu�o � s�N�� NN�_ì<:uJ�*rK���� rA�F �<;t��a t:�Q t4</t0<,u!�r�j� �! �<;t��< t�, t</t� N�ø ��N��P���C����&�CX�< t<t<
�< t<=t<	�PSW��2��&Ƈ &8u&� _[X�<r��SWV�����>�u�
�t��2�� &��
�t�^_[�SW���ٷ ��&��!_[�  �>Xcu��ar	��fw ��WÀ�Ar	��Fw��7À�0r	��9w��0���SQ�3�3�3�3��Xc
 &���r0
�u&�L��xt��Xu�Xc FF&�F��r� r��r����N�Y[�P���&Xcr��X���&Xc���3��X�Q��蒱���Y�V�R�!&�� =��t���^�P&� = t=	 t�&� =SCX�QR�����r/��3Ɍ�;�s(���uA&�  <Zt��& @������& ;�s3�I��ZYÃ>Xcu	��=��u@�PS�Y�� X�!��&�B% P� ��[
ظX�![X����<�u���
�t���PQ�r9������&��) <�t 3�A��s���� r����� 
�u�
YX�����SV���2�!��Ë�^[�SV��2�!��Ë�^[���&��R������t���Z�P�| r!��t�* u�, &�  <Zt��& @����X�P���
�X�&�  �&�  &� HI&�
 DD&� EN&�   �P&�   �  &� &�
 &� &� X�PQR2������3�;�t��uA&�  <Zt��& @�����ZYX�SQ���r93�3����t'�t�u&; ��&� &�  <Zt��& @���ԎË��u�Y[�P2�������
�X�SQ�،�&� �� ;�wE&�  &� &� &�  M�@����+�H&�  &�   &� �  &� &�
 &� &� ���Y[�SR����t+���>�r$P���M�[�t;�v��������t	�t�r���	���V�u3Ҋ��X��t����Z[�P���r��� u��&�  <Zt��& @����X�P&� = u"&� =FRu&�
 =OZu&� =ENu&� =  X�&�  &� FR&�
 OZ&� EN&�   �PQR�o�2���Z���3��k�uA;�t���u��&�  <Zt��& @����ZYX�PS���
 ����[X�PS�R�!&�G���&�  <Zt��& C�����=��[X�2����A�X�!2����B�X�!�� r�u � r���M��Ǿ� �����s= u����ú��= t������ ÿ-��  �<*t(<?t$<t:	�t
�t< t
�t�A��2���tN�ú���ú���ÿ� 2��ɬ���
�t<u�&�� ��#��%��%�á��H� �����C���IPQ�ȿէ���������- YX���c��t= |�ú���� �����������.>I&T_}�������#�:�L�]�y��������������9 at����	�
��#\m}�����6Y c!n#w$x%x'�(�)�*�+�,�-�.�/�0�1�2�3�4�5�6�7�8�9�:�;�<�B
CDE(F9GRHkI�J�K�L�M�N		O?	PV	QV	�W	T	(�	)
<�
=�
>7P�x�yvz�{N|�}�~j��-��������o���A�\�����z�������C�������w������s�G��M~� ,f@�A�BT�UV�h�i�|t���������.����N 	� � 0!0�!D�!EU"F�"G#H�#I$J{$X�$YS%Z�%[ &l�&��&��&��'�L(��(�J)��)�*%1 bytes free
#File cannot be copied onto itself
Insufficient disk space
Invalid code page
Invalid date
Invalid time
Invalid path
!Press any key to continue . . .
Unable to create directory
!Volume in drive %1 has no label
Volume in drive %1 is %2
Volume Serial Number is %1-%2
'Duplicate file name or file not found
Invalid path or file name
Out of environment space
File creation error
Batch file missing

Insert disk with batch file
Bad command or file name
Access denied 
)Content of destination lost before copy
$Invalid filename or file not found
%1 file(s) copied
%1 file(s) Invalid drive specification
&Code page %1 not prepared for system
+Code page %1 not prepared for all devices
Active code page: %1
NLSFUNC not installed
 Current drive is no longer validLabel not found
Syntax error
Current date is %1 %2
SunMonTueWedThuFriSatEnter new date (%1): Current time is %1
Enter new time: ,    Delete (Y/N)?<All files in directory will be deleted!
Are you sure (Y/N)?MS-DOS Version %1.%2Invalid directory
6Invalid path, not directory,
or directory not empty
Must specify ON or OFF
Directory of %1
	No Path
Invalid drive in search path
Invalid device
FOR cannot be nested
%Intermediate file error during pipe
&Cannot do binary reads from a device
BREAK is %1
VERIFY is %1
ECHO is %1
off on Error writing to device
%1%1%1%1	
 <DIR>     
%1	mm-dd-yy 	dd-mm-yy 	yy-mm-dd %1 %2%1 %1  %2Directory already exists

%1 bytes
Total files listed:
*(Error occurred in environment variable)
 [Y/N]?YN(continuing %1)Revision %1
DOS is in ROMDOS is in HMADOS is in low memoryCannot Loadhigh batch file
LoadHigh: Invalid filename
0Cannot open specified country information file
LoadHigh: Invalid argument
Required parameter missing
Unrecognized switch
%A bad UMB number has been specified
  %1.%2 to 1.09                 %1.%2 to 1.0 average compression ratio
Overwrite %1 (Yes/No/All)?YNA     �Sets or clears extended CTRL+C checking.

BREAK [ON | OFF]

Type BREAK without a parameter to display the current BREAK setting.
?Displays or sets the active code page number.

CHCP [nnn]

p  nnn   Specifies a code page number.

Type CHCP without a parameter to display the active code page number.
[Displays the name of or changes the current directory.

CHDIR [drive:][path]
CHDIR[..]
bCD [drive:][path]
CD[..]

  ..   Specifies that you want to change to the parent directory.

�Type CD drive: to display the current directory in the specified drive.
Type CD without parameters to display the current drive and directory.
Clears the screen.

CLS
�Copies one or more files to another location.

COPY [/A | /B] source [/A | /B] [+ source [/A | /B] [+ ...]] [destination
  [/A | /B]] [/V] [/Y | /-Y]

h  source       Specifies the file or files to be copied.
  /A           Indicates an ASCII text file.
v  /B           Indicates a binary file.
  destination  Specifies the directory and/or filename for the new file(s).
?  /V           Verifies that new files are written correctly.
t  /Y           Suppresses prompting to confirm you want to overwrite an
               existing destination file.
r  /-Y          Causes prompting to confirm you want to overwrite an
               existing destination file.

BThe switch /Y may be preset in the COPYCMD environment variable.
�To append files, specify a single file for destination, but multiple files
for source (using wildcards or file1+file2+file3 format).
�Changes the terminal device used to control your system.

CTTY device

  device   The terminal device you want to use, such as COM1.
]Displays or sets the date.

DATE [mm-dd-yy]

  mm-dd-yy    Sets the date you specify.

�Type DATE without parameters to display the current date setting and
a prompt for a new one.  Press ENTER to keep the same date.
dDeletes one or more files.

DEL [drive:][path]filename [/P]
ERASE [drive:][path]filename [/P]

�  [drive:][path]filename  Specifies the file(s) to delete.  Specify multiple
                          files by using wildcards.
O  /P                      Prompts for confirmation before deleting each file.
�Displays a list of files and subdirectories in a directory.

DIR [drive:][path][filename] [/P] [/W] [/A[[:]attribs]] [/O[[:]sortord]]
    [/S] [/B] [/L] [/C[H]]

P  [drive:][path][filename]   Specifies drive, directory, and/or files to list.
Y  /P      Pauses after each screenful of information.
  /W      Uses wide list format.
~  /A      Displays files with specified attributes.
  attribs   D  Directories   R  Read-only files         H  Hidden files
{            S  System files  A  Files ready to archive  -  Prefix meaning "not"
  /O      List by files in sorted order.
�  sortord   N  By name (alphabetic)       S  By size (smallest first)
            E  By extension (alphabetic)  D  By date & time (earliest first)
F            G  Group directories first    -  Prefix to reverse order
            C  By compression ratio (smallest first)
  /S      Displays files in specified directory and all subdirectories.
A  /B      Uses bare format (no heading information or summary).
  /L      Uses lowercase.
R  /C[H]   Displays file compression ratio; /CH uses host allocation unit size.

�Switches may be preset in the DIRCMD environment variable.  Override
preset switches by prefixing any switch with - (hyphen)--for example, /-W.
    [/S] [/B] [/L]

  /L      Uses lowercase.

>Quits the COMMAND.COM program (command interpreter).

EXIT
=Creates a directory.

MKDIR [drive:]path
MD [drive:]path
]Displays or sets a search path for executable files.

PATH [[drive:]path[;...]]
PATH ;

kType PATH ; to clear all search-path settings and direct MS-DOS to search
only in the current directory.
;Type PATH without parameters to display the current path.
7Changes the MS-DOS command prompt.

PROMPT [text]

|  text    Specifies a new command prompt.

Prompt can be made up of normal characters and the following special codes:

/  $Q   = (equal sign)
  $$   $ (dollar sign)
*  $T   Current time
  $D   Current date
=  $P   Current drive and path
  $V   MS-DOS version number
4  $N   Current drive
  $G   > (greater-than sign)
,  $L   < (less-than sign)
  $B   | (pipe)
y  $H   Backspace (erases previous character)
  $E   Escape code (ASCII code 27)
  $_   Carriage return and linefeed

LType PROMPT without parameters to reset the prompt to the default setting.
GRemoves (deletes) a directory.

RMDIR [drive:]path
RD [drive:]path
Renames a file or files.

SRENAME [drive:][path]filename1 filename2
REN [drive:][path]filename1 filename2

�Note that you cannot specify a new drive or path for your destination file.

Use MOVE to rename a directory, or to move files from one directory to another.
WDisplays, sets, or removes MS-DOS environment variables.

SET [variable=[string]]

�  variable  Specifies the environment-variable name.
  string    Specifies a series of characters to assign to the variable.

KType SET without parameters to display the current environment variables.
-Displays or sets the time.

TIME [time]

�Type TIME without parameters to display the current time setting and
a prompt for a new one.  Press ENTER to keep the same time.
FDisplays the contents of a text file.

TYPE [drive:][path]filename
%Displays the MS-DOS version.

VER
�Tells MS-DOS whether to verify that your files are written correctly to a
disk.

VERIFY [ON | OFF]

Type VERIFY without a parameter to display the current VERIFY setting.
RDisplays the disk volume label and serial number, if they exist.

VOL [drive:]
[Calls one batch program from another.

CALL [drive:][path]filename [batch-parameters]

r  batch-parameters   Specifies any command-line information required by the
                     batch program.
LRecords comments (remarks) in a batch file or CONFIG.SYS.

REM [comment]
kSuspends processing of a batch program and displays the message "Press any
key to continue...."

PAUSE
MDisplays messages, or turns command-echoing on or off.

  ECHO [ON | OFF]
W  ECHO [message]

Type ECHO without parameters to display the current echo setting.
GDirects MS-DOS to a labelled line in a batch program.

GOTO label

�  label   Specifies a text string used in the batch program as a label.

You type a label on a line by itself, beginning with a colon.
JChanges the position of replaceable parameters in a batch file.

SHIFT
ZPerforms conditional processing in batch programs.

IF [NOT] ERRORLEVEL number command
FIF [NOT] string1==string2 command
IF [NOT] EXIST filename command

}  NOT               Specifies that MS-DOS should carry out the command only
                    if the condition is false.
�  ERRORLEVEL number Specifies a true condition if the last program run returned
                    an exit code equal to or greater than the number specified.
f  command           Specifies the command to carry out if the condition is
                    met.
j  string1==string2  Specifies a true condition if the specified text strings
                    match.
g  EXIST filename    Specifies a true condition if the specified filename
                    exists.
wRuns a specified command for each file in a set of files.

FOR %variable IN (set) DO command [command-parameters]

}  %variable  Specifies a replaceable parameter.
  (set)      Specifies a set of one or more files.  Wildcards may be used.
V  command    Specifies the command to carry out for each file.
  command-parameters
�             Specifies parameters or switches for the specified command.

To use the FOR command in a batch program, specify %%variable instead of
%variable.
Reserved command name
/Loads a program into the upper memory area.

�LOADHIGH [drive:][path]filename [parameters]
LOADHIGH [/L:region1[,minsize1][;region2[,minsize2]...] [/S]]
         [drive:][path]filename [parameters]

�/L:region1[,minsize1][;region2[,minsize2]]...
            Specifies the region(s) of memory into which to load
            the program.  Region1 specifies the number of the first
�            memory region; minsize1 specifies the minimum size, if
            any, for region1.  Region2 and minsize2 specify the
            number and minimum size of the second region, if any.
            You can specify as many regions as you want.

�/S          Shrinks a UMB to its minimum size while the program
            is loading.  /S is normally used only by MemMaker.

W[drive:][path]filename
            Specifies the location and name of the program.

Zparameters  Specifies any command-line information required by
            the program.
�>0i��k-�     & ��6 File not foundPath not foundInsufficient memoryExtended Error %1�>����^��� Parse Error %1�>�����     %�   �  � � � � � � � � � � � � � '�  �		 � *�  �		 � .�  �   � � ��  � � ��  �   ��  �         ��        4

 	 
            �     2�  �  4�  �0 8�   �  8�   �  o�  �  ��  �0 ��  �0     >�  �             �       � !     � # $ % & ' ��  �  ( ��  �  ) !�  � * %�  �   + , Q - . 0 1 2 3 ��        4
 4     � 5     �
      � 6 7 3�  � 8 9 : ; < >�  �  B 6�    C D E F G H I J K L M ,�  �  -�   N ,�  �  -�   PATH=PROMPT=COMSPEC=DIRCMD=  ()  <=>  P  xyz{|}~  �  ��  ���  �������������  �  �       ,  @AB  TUV  hi  |  �  �  �  ��  �  �  	    0  DEFGHIJ  XYZ[  l  ��������  [2JBE$D >E9$G=$H/$LA$NV$P`$Q5$To6V�#_a,$G$ NOT�
ERRORLEVEL�EXIST  DIRg1�CALL��CHCP�&��RENAME� u�REN� u�ERASE )�DEL )�TYPE7!��REM��COPYm>�PAUSE���DATEn5#�TIME�5��VERa#��VOLe"��CD!+�CHDIR!+�MD�+Q�MKDIR�+Q�RD ,q�RMDIR ,q�BREAKf=��VERIFY�=��SET�(}�PROMPTg(]�PATH�$U�EXIT �'M�CTTY&�ECHO,=��GOTO5��SHIFT���IFi��FOR�ɚCLS u%	�TRUENAMEA'ӚLOADHIGH?hךLH?hך .COM.EXE.BAT-Y?VBAPWRHSvDANEDSGC        u�ʜ  u�ʜ  u�ʜ    u�ʜ/P ��  ��    u��    �f�ON OFF �   �  �  u�)� d   �    9�  ?�    }�ʜ K�  Q�    ��ʜ ]�  c�   ��ʜ o� ͜  x�  ֜  �� ͜� ��  ߜ����  ! u�̜/A /O /C     u�ʜ/-A /-O /S /-S /B /-B /W /-W /P /-P /L /-L /-C ܝ��ʝǝѝΝ����Ý��؝՝��������� ͜͜  � �     u�ʜ  �   &�    u�ʜ/R 5� ͜  TEMP= COPYCMD=\DBLSPACE.                                                                                                                                                              ��                                        �    �    []|<>+=;"             ����        ����        ��������            ����       
     
 $$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$MS DOS Version 6 (C)Copyright 1981-1994 Microsoft Corp Licensed Material - Property of Microsoft All rights reserved                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              MZ� �       ��    �μ�  @                                    �                                                                                                                                                                                                                                                                                                                                                                                                                                                                  ����Bh=�DBLSPAC,.�Uw  �=  �  ��  �|�  �cB  �B  ��  MSFT      �    �      $$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$.�B .�B .�B .�B �>  .�B  .�> .�@ �   .��  .�>�.���� �� r��� s��'��  v�  QW�����_��.�>�.��Z�ʃ����.��.����v��� .�&� ��X�����2��| �.�6.��� ����r$�� �C3��.�� u�!r
�=�!��r��� t��
�u�f
�t� ��
�u|�
�uu�
�un���>�!�� u��C� �!.�>�  u���� �� u�Y��A�U�J� �/�>X u���t��X�U.�� �P��>�!X���".�	�=:\u-�
� � � �
�
�t<.t�������� �����øD�	��@�!��t�Ȣ��                                                                                                                    C                                                                           MDA�                                                                                                                                                        �                    X:\DRVSPACE.000DRVSPACE000SQRVWU�v>�� ��>&�6R ���&GA�	�&�G��2�CA�FA��u#�EA2��DA,B���9��Au�^t	H�����6A�Y��
�t������d���������d�������;r���r����
� ���	�t&�]��&�]����t�� �Z���ãZ ��+�)��� �Z�)��
�u���� �.�N
�u��
�u��>

�us��� ����Z�������d�����>u�� �Y*DA2��U�~-�>X u.�Y��AR�Z
�u���>u
�	��A��Y*DA����v> ]_^ZY[���Z�?�> ��PS��>&�_�X���&�GC @[X��%r<��3���>��?���>��>������>;�>r��>������ @��  �����A�����G�G  �d�h��A% �� tH�3����������� 
��t��j��t��2��	��A�uv&�G��&�G	��&�G������&�G����&�G��&�GH��&�G��&�G��&�G��&�_���t#&�G��$��&�G�d�f&�G�h�j�À>v>u$��&�G&�W��� ���  �6����� B3�3ҋ�!�?�@ ��!� 
�t� �9H�& �����(3��t�5�7�>v>u	������B3�3ҋ�!P��3��6 ��X�6 - �� +@�� +<�� �\�^�S�3��6 ��3��6 ���@ ��&�l ��&�n ��2�áH.�� ��� ��u�>HtH��> t-= t;�>v>ti��� ��u\=  u�>v>tP��> u��C.�>� u.��  ��>v>t�"� ;�r= t���"2����u
=  t= t�ðÃ># t��>%u�>& t�>& u߀>*�u؃>+ tѡ13uȡ57�(t�u�@�t�2��MSDSP6.0MSDBL6.0�>� w>��3��6��ȡ�PQ��� 3��r#�>���WQ�
� �Y_t�� ��YX@��3��YX��YX&�E�����- ��2������ á\+��`�^��bs�\���^���`  �b  2����  ��  � 3����>�3����Q� ����� ��Y���������>� t� �� H��#��������;�r� ��R�������Q�����vY��Y�	���g3�����@���������������u= s� �>� u"������Q���Y��  �uj;�sf� �� J��#£��裯����;�r���6�������� �᣻�6��>�3ۋӡ������艷��������B����5�7�"2�;�s���H3ҹ - �� ;�s���@��3�VQ� ���� ��  �� �ʋ��&� ���I� ���u.�B +���𭒭��� �tQV�  ^Y��Y^F�3�.��Q�OY����2�Ëڱ���CP.�"2�.�.�� X��.+@�� rd- �� r\.+<�� rRPR.+\.^ZXsB������������������.;�s(.�6���PSQR�' ZY[X����uB.;�r3�@Ku��.��.�� �QR�- XY�ظ ���&�t.��.�� �.��.�� &	�.��.;��th.��I�$������.;�s�.;��tF���.;�r3�P�= X.���S.�&�. �� �ʋ��[S.���.���.������[��ğ��S����&� �� �ʋ��u��[S���;�ru������������[á �l�"2�n�b���9�p� 3��6 �r� 3��6 �t�#�v�<�x�>�z�@�|�B�~�D���;�������*����	,A���&�G���
��&�G�
,Т����R�������$ �������� �����t3Ҹ��� ����J� �/�u
;�s����������Z  ���M��&�G&�W��2�&���� ��H;�u���&�? �r1�����;�v�	 á�������&�G&�W&�  ���2�&����= r���+��� s� Á>����r���9�s�r���- � ��Z3�Á>��s7������3��; �6�&� C;�uP��@�3 X�6�&�$�s���%��3���� � �6�&� ��6�R�� [�;�t��3ҹ ��� À>v>t"�����������	,A������%X��p>��?����?��>��>�N'���<ar<zw$��3��tA��s�I���FAT16   �%�+5�7 @>���-���/�<�& �ʋ�QR��R,�$2��� �����$ ��>�� ���>���6��Ȏ���.�6��t'����� �2��ZY�4� ���`�<@�& �ʋ�QR�� ���7�>�����&�=DRu.�����>� t����ZY�� � ���2��ZY�ù 3�������r.��&�G��&�G��&�G��&�G'��&�G)���>v>t�&�G��&�G��&�G������&�G��&�G&�O2���&G�����H3��6����P2���[���X&� t
&+G�����V&�w &�W"+��� �t��������^���À>v>u��PR2������������ZXø B��!ø ?.�p>�� @.�>� uN.�p>.�>v>u9.��>��>������ȋ.���- �� ��� ��$�Āt���.��!�                                   ��������������������������                                  �  P��>&�R ����ğ�&�G����&�G������>&�R ���&�N &G2䓀� �t&�g��t��ty��tg��tX.��.�.�� �`t�>�?�tS�ذ����[<�t�&�GX��� &�G< "&�g��>&�R ����
�x����u���X[��t�&�G X�� u�� �� ��r��> &�G&�_�� ��&�`ul�� ug� QRVWUS&�g��A�������3��&�G�������A��r	�>�A�t�[]_^ZYr���o �r&�G����=����������&�G�<X.��.��SP��>&�N �<&�G�&����;u��?�&�?����Ћ&?��&����;y
���?�&�?��&�S2���;��A[��63�65#7#9�3�5SV�� �2����� �C��^[YZ� 
 Pe{����Lg~�
Cannot run SMARTDrive 4.0 with DriveSpace.
$�uO����tIPS�Ќ�;�u�>q��u�>� [Xu-�t�	�!� L�!�.�> A t���.��>�3 ��π�Jt=t,=t=�    <t�<t�<t�<u��!��� s/�.��\���u.�z>�.��v&�P3�.�z>.��>.��>X��3��MD.�Z.�DA.�.EAϸ��s��2��.���A3��3�.�>{>t��!��� �P��!X�.�{>�J� �/.�{> Ê�2��.���A�Àt��W����.:��At��_����S���r%.*DA��A.:EAs�.���>�MN�E�u
�}[ϱ���
�uPS��r�.*DA��A.:EAs�.8�?u.�6?.�?.�>?.�?.�T?�.���>�w
�G��G�WN[ϸ��sN��2��.���A�ƀ �t:���.���A:�t	�;Ƹu#.���A$�
�.���A.���A�Ɗ����� ����&�|Au0��2��.:��Au#��.*DA��A.:EAs�]2�RV�(^Z�]�&�D��E�i�Iϊ�� �t�2��.���A�t6.���A% �����.:��Au��.*DA��A�6?.8�?t��.���>3�ø�.��>.��>3��U�>~>�>�>Zp>����Y�ʋ�.�.9B.�CA3��.�>w> t��3��3�3���.�>w> t�.�3.�5��.�&B.�&0B�B� 
�u�'B�
 
�u�& 2�ÊT	�N �u�\�D&�G�D&�_��D2����>!B�'B� �>+B�B� �ÊD&�E&�E��&�E�D&�E�.��>&�&:t��&�?�u���S.��>&���S.��>&��.�>�>�uP��QR.��>ZYX[� �.�>4A ujWP3��ǿh &�E&X_t�P���X��CIuԁ�MRu�&�E �t�.�4AV�"A��� �^&�e�&�E.�3 &�E
.�5 &�E2 &�M
��"A�CI�MR� S&�^ 2��.���A�u[�PW.���A% �����.:��Au��.*DA��A�>?.8�?t��.���>.�} t�_X[�.�}� w�3����                                                                                      
              �<D[W��	����@A S�܀�lwY2���T���
�uK[�ڊg��S�ܴ]��]t5��<u/�5A [VW����t�
�t��u.�5A_^�[�.�.J�t>u��At��� ��
�t�[��.�J�.�t>u.��At� �U��r�f�]πN]�Z� ���w���
[U��]t�R��.�J=��tۋ�[VWPR��riP�G��Xuk�؋T�D�u=� w3�;�s!��Q�DF�TH�|�L��Y�t�������������ܻ���	��;�s����;�vZ+�����ZX_^]��P��g ��X댋���PSQRVW3ۋˊDA��A��ۊEA���A�u;��AuCCB����#���A�����9A??�D�
 �6A� �>9AKOt�_^ZY[X�.�R��U��P���&�� �F��&�� �FX�]��.�JU�윏F].�R�&�� &�� ��.�@A.�.N��t�&�}� t�&�}���V�  �ވ  P�&  �����u.�  U��f�V�  �ވ  �  �  P�&  ��Xu� ���.��?u�.��?.��?�aw�*(#]


]]

(#UUE


3 


���PSQRWVU�.��?.�&�?��Ȏ�.�&?�.��?�G.:EAsY.�&�?���t(.�>�? t �u:�tP�.��?X:�u.�x>�5�G�<w�W����G.��?3�.�>5A u.��OX��.��?���G�>x> te��?&�uZ�y>���uQ&�_&�G uF�p>��>��?�>�>3���>����>��?�Q�Āt��?&�G�x> ���?&��6�>�7?���9B@t�?�?4t��k���?�&�?�]^_ZY[X��?�>x> u��x> ��?&�wP.�T?&�GX.�?.�?.��?&�GˈG��Luk�.�>]?u	.��? �
�t
x.�>Z? u�G3��.��?�Gp?�O�����u-.�Z? .��> �G�O3����u.�>]?t� ��� ����u�9Gt��t.8�?u�.��>  �G=��u
�G.��>�G.��>R.��>.��>G�� - �� .+L?.N?Zr	�^���Q�.�>�> u.��>.;(?r�)�w�W��Ɏ�u���.��?  .��>G.;(?v.+(?.��?)G�G.�p>.��>.+:?s��;Gr�G��.��>�� u� .��>.+:?.+B?s3�؋O;�r��.�>p>t.��>Q��.�p>Q��Y.�p>Y.��>� tZ.��>.+:?.+B?.+B?s6�؋O;�v��.�>p>t.�>.�7?��G)Ot�.��>.+B?�< t.��>.+B?�O�+ .�>�? t.��?�G.�(?.��>.��>  ���.��?�G3��)O.$?H+�W.��>�W.��>QS��[Y.�>.�7?��G� �� u���O.:�?u3��SQ+ۊ���.���>�Q�[X.��?� [��Y[����VWQ��?�> ��Y_^�G&��>�?H��>�?�S?�࣒>3���>��A��A��A��S��A��T?��G�G  �V?�G�?�?��A�Āu��A
�u�� u	�P u2���� [�����p>��>��?�>�>��?��>  ��>  ��Āu�&�E'9^?u&�E)9`?�S��>��>��>��>� �p>�$?3����>&�?�Du&�Ru�l?&;Gu�n?&;G[�.��?2�.DA��A.�y>S�.���A�u.�y>R��Z���� Z3���>��A�r>�q>���H�u&�G ��	.��?���t=*���.���>�t0.�?.�G.�?.�G.�Z?.�GT.�h?.�Gb.�j?.�Gd.��?.�Gz��	.��>  .�p>.��>.��>.�6�>.�6�>� 3�.�$?- �� ����'��� �����3������V��^�|?���p?� �2���Ȏؾp?��?2�ۋ��>�}j� �.�p>� 3�.�$?- �� �&3�Àu�ft��Ft��`t�gt����_C�+���_��G�G  �G �G���.�6�>��� .��FC��+���w&�<MDt� &�D<Fu�d�u<Iu6�Ȏ��W��>  �����k?�3۹ ���>�t���Ge��ڃ����;<Su=�_�Ȏ�2����㋿�>�t(�U&�T&�\�Ub&�T	&�\�Ee�t���J&�DKO3�É6�A��A��A��>+B?��A��>  ��A�>�A 3�á�A��A�6?��;�>u�>�At��A;�>t���X��A ��A �>�A t���A  ��A ��A ��A��A��A��>����>��A�.�>�.�A�� �u@�� u�t*�>�? u#�6�>UP��A �g��AX]��>��>�>u�X��A  �"���?��>9�A}� ��At� ��>�A t'���A�6�A���6�A�>u>u���7r>�>�A�?)�A��>  �A��A +�Av�Q?������3��>�A��A��>�A��3���A��>��A����������؎��6�A��>�A t�>u>u��A�6�A�r���=��A��A#�>�;�A|��A�>u>u��A�| �>�A;>�Aw�>�A�?+�t�Q?��������>�A�3���6�A#6�>��A�?+�;���)�A�A��A �>�A��A�Q?����6�A������>�A����A���;�|�9�A|P�%�ʋ�A+ˁðA��A�? u� ��r,�� C��ځðA+�uÀ? u�� ��r	��ACHu������ځðA�? u�CB;�At�;�|��SQVW��A�7�>�A#>�>;�}>�A;�|+>�A�����A�  �? u��@SQR�M�ZY[CB��_^Y[�PV�؎��6�>��^X�P��A��A��AX�PQW�Ɏ���>��>�A3���_YXá�>+B?��A��>  ��A��A�k?�t��
�>�A ~0��A��A�6?��;�>u �>�Au��A;�>t
��>��>��>�� 3����A ��A �>�A t�5��A ��A �I���>���>��A��>��A���A  �>�A#>�>uR��A;?|H��>%����@��A�?��A��A��A��A�6�A�?)�A�A��A 6�>�>�A u�� �� ��>���3��>�>���>�.�>��A  �� �t*��>u>u���>�A tV�6�A��^s�����]��A �>�A u�*���A�6�>��A��A�>�A#>�>u��A;?|�����A�?+�;�A~��A)�A�A��A ���;�Ar��A�߁ðA���C���Q?����>�>���،Ȏ��������>�A u�j?h?t�6���A V�
 ^��A�"���A;�A��A��A��A�6�A�ȡ�A��>��A��>��t3��A �>�Au;?u��t��A����.�>�A�u> �>s>u�s>�Q?����A��u>�؎��6�>�F��A  ��A ��A�.�A�� �u<�>@A tU�� u�tK�s��AH�Q?��@;�?u7������>�? u'���^�d�6�A��AH�Q?��@;�tQ��>��>����6�A����u?��> �t�6�A��>��>����>�A t� ��>  ��A ���'����.�>��>���� ��6�AN�Q?��F�6�AN����6�AN�
���>s> t�� @��>�.�>��A�.�A��A��A��>����A���p>�6�>��>�6�>��>�>s> t��>�+3����A �8���A��6�>��6�A��>S��>P��%����@��A��X�p>��>�6�>�; [&�?JMuP��% <�
��@��AX�[�&�?DSt���A  ��>  �>�A t�������u> �� @t�u>S��>&�JM&�G  ����>[U���{
]�PQV�* �I^YX�.�6�?.��?�+.�&�>����.��?��.�&�>��.��A PQV.�>�A tSR�Ȏ��E�Z[.��A".��A-.�>]? t��.�>t> t	.�p>�0^YXÀ>�A u��>  �PSVWU�>�A t����>  ��A ��>�.�>��A����A r<�>�A t5���6�A�>�A;>?s�Q?��>�A� ������3����j�6�A�]_^[X� QVW�ȋ6�A��>�>�>�����A��_^Y�P3�� ��A��AX�S��A��G�G�G�G�G
�G�G[�QVW��>��ΎƋ6�>���>�>��>������?��A��A_^Y�P�@ ��&�n .;�Awr&�l .;�Ar.��A &�l 8.��A&�n   .��AX�PSQRW����A�?&�= t\&�}  tU�>�At�? t>&�} uB&�}L u;&���  u3&���  u+&�� u#&��L u&��� u&��� uC>?���3�_ZY[X�.�9B tVQP� .�6~>.��>�.�1BXY^�.�9B t9VQP.�>r>�t+� .�6~>.��>�.;1Bt@���u.1Bt���XY^�.�9B u��5�O.1B.�1B 5�O&�5�O.)1B.�1B �.�9B0 tVQP� .�6�>.��>�&.�3BXY^�.�9B t1VQP� .�6�>.��>� .;3Bt@���u.3Bt��cXY^�.�9B  u�Á��O.3B.�3B ���O&����O.)3B.�3B �.�9B tVQ&�&�u\��+�� Y^&�E`�.�9B t3VQP.�?��.�6b?+��p .;f?t@���u.f?t���XY^�.�7Bu�.�7B
 .�Z �u�.�9B t1VQP�p>�Z+΃��� .;5Bt@���u.5Bt��XY^��SRW��O3�3����� t�3���I�� u�����t�3��ڭ3��ڭ3��ڭ3������_Z[� @��?u3ҋ��P�>�?t�r>��:P?r*��r
X�+PSQV��>���>r>�u*��W
����P?��?N�Q?��F��? 2�r>�&�/��и �3��~>&�?��u3�����;�>r��x����� &�t3���s���G;�u�;.
?wr;?r��?�J�)6?�? +փ� ��? &�?��? P&�t�X��s��Nu���� (?�� +B?�� $?�� �q>�k?�uR��?��h?j?Z���^Y[X�PSQV� r�6?�? ����? P��&#��X&�?��? ��r��Nu��PSQV�] r�)6?�? ��? &�?��? ��&�����s��Nu��m�PSQV��?�" r;�>s&�u��s��Nu���? ^Y[XÎ�>�M �5�+(?�� B?�� +$?�� - �� ;
?w'r;?s�6�/��ڱ����~>�ʀ�� �������P��?:�?t��?�r>�X�SQVW��>������]�?�
?�6�/�t����?3�3�2�R�?Z��>~>� �>�?u`R2��&�/�6?+��Ƌ6
?�ֹ ���t;PS���ظ &�u)&���>�? uW�6�?��?�2�&�>�q>�2��?_[X��Z�3������+�ރ� �u�r>����?t�i��ãh?�j?�r>�P��X_^Y[�.�&�>��>�q> 린����	&�D�*_^&�D�..�;BQRVW�j�r�.�;B&�D ����.���> u�&�D3ҹ ��@.;�>w�+�.�CA�FA.�|>.�=t
| G��u��.���>.��WA.��WA1.���FA�߃����ٌɎ����| ���&�Ee�SW&�� �P3���.��>.+�>.)�>����&�u\.�>�>���Y����_&�E\&.��>&�E^[&�]V.�\?��S�_R2�ۊ��A[�GR�gS�P����j�X.�;B.DA��A���.���A�� �ڸ �8.��?�.��?�_^ZY3��P��>&�_�X���X��% @&�gC��&	GCÊ�2�ۋ��A�ǀ t1���8��At&R2���Z�ڸ �� *DA��A��2����.���> u��S2��.DA,A���.���A���r�{���[r�.Ǉ�>  .�\?*�.ƇFA.��?�.��?��?+b?� ���3����>��>;�>vT+�>P�b?+�>3���Z+�t?����6?�>b?�ȡ�>�؎������ ��3ۋb?���>�t
9U\v))E\CC��3��.�>z>uP.��>.�>tX.��>�SW3��Ǹ��; �/.�>�>.��>���_[Xt��� S�V��6b?+�+��	;6?w4��&�� ;�r�w;�v�&++�&�D��>&�D��>�>��> �[��[�SRVWU�ʎڋ>�>�>�?�>�> �� �يU?*��������������r2&�+�Q�?�U?��Y;�w2��?�r � �u3�]_^Z[�.��?���.�&�?�.��>  ���?�@ � �u�+˃�;6?w�&�D��>&�D��>���u�&��.�6�?.��?N6�D�.��?��SQRVW��?.��A.�>�A.��A�T?.��A�p>.��A.��A  �V?.��A��?2�.��A�>W? t.��A��.��A��>.��A��>.��A���>.��A��A�?�?��A_^ZY[�SQR�ӱ	��:�?t�>t> t�p>����?�p>������	��+������>��>&���>&�O��߉�>ZY[�PSQR�ӱ	��:�?t�>t> t�p>�u��?�p>�i����	��+ڋ�2������>��>��>&9t�������>���&9Ot���������
�t�ڊQ?����Ƈ�?�t>ZY[X�PS.��?�G<t<t<	u�G  [X�PSRVU�.+"?.�>[?u�|.�Q?�������.�*?،ʎ��Nr+&�= u(���.�>��>�� �t���&�>������C���.�>@A t����.�>��>�� �u��� u�t�;�>t����Z�� R.�&?��.;�?s�.�6�?�t@=�s܋�.���?.��?��.��?ZP��.�&?��.;�?r���.�6�?��X��+�;�s��.�*?،ʎډ�?�| s�q&��>�? t���%�u1����.�>��>�� �t� �� �&�>����6�?uGGC��?t/�.�>@A t����.�>��>�� �u��� u�t�;�>t��4 ��]^Z[X�.;*?r"PR.�?��.B?�� .+L?.N?�ZXr�:���Q�> �6�?���|��>�? u$��> @u���r�>�A t���&���> ��r�Y�3���>��>��PQ��%����@��?YX���Q�6�?��.;�>u.��>  .��A ��Y���?��t> ��?  ��?  �PQU:r>tJ�>q> t�D �>t> t�p>� �q> �r><�t%�& ?+��p>��>��>�6~>��>� ?�.����]YX�.�>q> tN�J�PSQRU.�>r>�u� �$.�r>.�& ?+�.�p>.��>.��>.�6~>.��>.� ?���.�q> ]ZY[X�PSQRU.��>.��>.��>.��>.�?3�.��?��.?+�.�>p>t2�V�.�?��?.�?t
I.�>@C��?.?.�?tIK���m��.�6�?.��?��]�X.��?��.��?  .��?  .�t> ]ZY[X�.��?.��?��?P.��A$A.��?��?&�G&�O��?&�G
&�O��?.��?.��?3�&�G&�GX�P�'=&��?&��?��?&��?&��?X�P�`.��?�a����a���a�� � �X�S3����&�$ &�& .��?.��?�<&�$ &�& �[�PS3���.��?.��?�&�$ &�& �.��? [X�.�F < t<
t<u�+ �� E��ôP�c X��Q� �	�W Yð ��P���X:�w�ôP�����2��P��������� X$�':'.�C�P�� �� .��?.�6�?X�.��?.�6�?���.�&�?SQRVWU��?��.��?]_^ZY[��/ ��3ҳ��?S�H����.�>�?Nu���[� ��?3��/���.��?�WSP3��ǻ ���/���t�z=PW� �X[_��PSQR� �@ ��@�� t�s>�>AZY[X���s> �6�@��@�Q?���@��>��@� A��>�A�P��>�P��A �
A�A�6A�A3��A�AX�PQ�ƊQ?�����>A�6
A����Ȏ؉6
A�>A�YXÀ>�At�PSQR�Q?��6A�AAu�.
A�A�
A� u�>A�>A t>A�ZY[X������@� &�_��                                               ��                                                                                             �u��                                                                                                                                ��        �  �         ]6                               C:\DRVSPACE.BIN                   DoubleGuard Alarm #00

A program has corrupted memory belonging to DriveSpace.
Further disk activity could result in the loss of some or all of the
data on your drive.  Therefore, DoubleGuard has halted your computer.
For more information, see the README.TXT file.                                              �                     MDF??12345                                                                                                          -                                                 �>                	 
                                          
     C:\DBLSPACE.BIN C:\DRVSPACE.MR1     �=Jt.�.^B.�> A t��RMu��ICu����.��>�< &�]ϝB  �� ˸ �S��.! A[�.�.�B@t�H.� At��.�>qu u�.��>�&8r��.�qu&�.�pu�.�&lu.�nu��ʎҼlu��" �.�nu.�&lu��.��>.�pu&�.�qu ��=  t=@ t=� t= t
� �� � �u  �B r7V�4�j�	� �vu��%�t���vu�/^;|s�|.�>ru u3�ø ø �ËD�t&�б	����|&�JM&�E  �T��Jr.�p����V�D�б	����t@.�su�|�4�3ɭ=JMu��.�zur^+|�|3��=DSt�^� �V�D�б	����t@.�su�T�\�|�4����u3�=JMu:��P.�zuXr3��^=DSu�΀�T�\��ǇD+��|3�øJM�ƀtθDS��=DSt��   �DE�E�EgF�FJG�G.��> tS.��>�Ã.�su.��>�[.��>���=DStғ�u�+�� �˽ � ��.��dD��u��Mx�������u<�u�б���?����5�u�б��2���ă�@���б������@�!�p��Mx��Ȫ���Ĩu�����$Mx᪬������uC�u�б���?������u�б��2���ă�@�%���Э�ȃ�ѱ�ʁ�@�������Mx��Ȫ����ƨu�����$Mxݪ�������uC�u�б���?����D� u�б��2���ă�@�%���Э�ȃ�ѱ�ʁ�@�&�
�����Mx��Ȫ����ƨu�����$Mxݪ�������uC� u�б���?������@u�б��2���ă�@�%���Э�ȃ�ѱ�ʁ�@��'
�����Mx��Ȫ����ƨu�����$Mxݪ������� uA�@u�б���?����O��u�б��2����@�% ��Э�ȃ�ѱ�ʁ�@�/�	�����Mx��Ȫ����ƨ u�����$Mxݪ�������@uJ��u�б���?�������u% ��Э�ȃ�ѱ	�ʃ�@��% ��Э�ȃ�ѱ	�ʁ�@��D	�����Mx��Ȫ����ƨ@u�����$Mxݪ������騀uK��u�б	���?����^��u% ��Э�ȃ�ѱ
�ʃ�@�u% ��Э�ȃ�?ѱ
�ʁ�@�0�������Mx��Ȫ����ƨ�u��$Mx᪬������uH��u�б
���?��C��u% ��Э�ȃ�ѱ�ʃ�@��% ��Э�ȃ�ѱ�ʁ�@��^��Mx��Ȫ�����t��?t�t��xދ΋�+�&�&�&�������+� ��ڨt&�б����ʃ�+�x��֋�+�����x����t#�б����ʃ�+�x�֋�+�����*��t1�б����ʃ�
+�x��֋�+���t������������t1�б�����ċʃ�+�x�֋�+���t�������������t���?t�t��x��΋�+�&�&�&����L��=�� �ڨt&�б����ʃ�+�x��֋�+���������t#�б����ʃ�+�x�֋�+�������t4�б�����ċʃ�
+�x��֋�+���t������������ t1�б�����ċʃ�+�x�֋�+���t��������������t���?t�t��x��΋�+�&�&�&�������L��/�ڨt&�б����ʃ�+�x��֋�+�����u���t#�б����ʃ�+�x�֋�+�����8�� t4�б�����ċʃ�
+�x��֋�+���t��������\���@t1�б�����ċʃ�+�x�֋�+���t��������������t���?t�t��x��΋�+�&�&�&����H��[��>�ڨt&�б����ʃ�+�x��֋�+��������*� t&�б�����ċʃ�+�x�֋�+�����A��@t4�б�����ċʃ�
+�x��֋�+���t��������������t1�б�����ċʃ�+�x�֋�+���t��������}������t���?t�t��x��΋�+�&�&�&�������g��J�ڨ t&�б����ʃ�+�x��֋�+�����}��6�@t&�б�����ċʃ�+�x�֋�+��������t4�б�����ċʃ�
+�x��֋�+���t��������R�����t1�б	�����ċʃ�+�x�֋�+���t�����������	����t���?t� t��x��΋�+�&�&�&����B��r�
�U�ڨ@t)�б�����ċʃ�+�x݋֋�+�������>��t&�б�����ċʃ�+�x�֋�+����� ���t4�б	�����ċʃ�
+�x��֋�+���t��������������t1�б
�����ċʃ�+�x�֋�+���t��������r��
����t���?t�@t��x��΋�+�&�&�&�������y��\�ڨ�t)�б�����ċʃ�+�x݋֋�+��������E��t&�б	�����ċʃ�+�x�֋�+��������t4�б
�����ċʃ�
+�x��֋�+���t��������;�����t1�б�����ċʃ�+�x�֋�+���t������������� ��t���?t ��t!��x��΋�+�&�&�&��������|��_����t)�б	�����ċʃ�+�x܋֋�+�����V��G��t&�б
�����ċʃ�+�x�֋�+��������t4�б�����ċʃ�
+�x��֋�+���t����������� ��t/�б�����ʃ�+�x�֋�+���t�������������Q��ـ������sX% "��+�xI�֋�+���t�������ZЀ�rF���ҷ ��.��dD��sN�����ҷ ��.��dDY�C��s
%? B�����s% � ��
���sܴ ��녅�u
.�sut
�<�.�suu����                 �>�o�.p�p��t	���s�Ī+>�o�PSQVW���p�p  ��o�6�o��o�>�o��o�� ��o�����t�����6�o���>�o�ru ��_^Y[X���>rut3PSQ���6�o�o�&p���. p��r&�&�T���Tu��T� �ˇۃ�r�&�&�T��T��o��o;th����];t[����];tN����];tA����];t4����];t'����];t����];t����];u�:Gu����ou2���ls�m�����������E�ֈu���T������lPFI�A��ֆw���T�����놗�l����+߁�?s�S�������ٌڎ�o��tNA+�S��S���r&�PIu��. p� �P��o�.p���>�o�.p�p����^ ��
�yXz����s%ۋ�*���ƀ�6&����̀���À��"��ۋ�*���Ɗ̀�	&�����À��^ ��
�x���@s)��ۀ���*���Ɗ̀�	p&�����À��a��@s.��@���ۀ���*���Ɗ̀�<&�����À��-��@���ۀ���*���Ɗ̀�&�����À��^ ���� w,��pۋ�,p��*����*�&��������À������?s*C���� ��*���Ɗ̀�&�����À�� ��s)C����@ ��*���Ɗ̀�&�����À��x��� s)C���󀀋�*���Ɗ̀�&�����À��I+ҋ�*���ƀ�&����̀����C�����*���Ɗ̀�&�����À���������*���Ɗ̀�&�����À��.p�p�>�o�&pY[��op;�orX��ru���QW����T��o&�&�E&�E&�E
��Iu�� p�T_Y��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               																          ( 8 H X h x  0 P p � � � � 0Pp������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          Q  �D  �T  �T  4
DRVSPACE.BIN cannot be loaded from your CONFIG.SYS file.$  DRVSPACE.BIN was unable to load.
$You pressed CTRL+F5 or CTRL+F8 to bypass DRVSPACE.BIN. Therefore, none of
your compressed drives are available.
$
You are loading the incorrect version of DRVSPACE.BIN for this
version of MS-DOS. Since this configuration is untested, you
should correct this problem as soon as possible. Press ENTER
to continue starting MS-DOS.
$              ��                  ��u����.;Zt= r=2 r���[v�� �<u��Ȏ؉�?��?��� �� �գ�>�  �  �k�4�!��>��>��?�W��A�DA�
�t����,s	��u�	�!�����tHtD�{�>\w t;�@��dD��P��dD�l���P��T��P�dD�tD��dD��-@�dD������9�T~�dD��P��dD�����P��T��P�dD�tD��dD��-T~dD�����>CAv�CA�FA�CA*��G���UA��u�� �|>�|>�G1� �WA�CA2�| ��|>� ���ãrչ$ �|>�&�8w��W��>&�D 2 &�F ��B��>�< �>�@��@_���ر���ȃ���>��>��>��>��>� �� ��裲>��> t�>� ��>�R�!��>��>�a 3��� ��u� .��?�G �G  �O.�   � � �?��>�( ��>�( �~> ��> ��> P��>��A��>��AX�R.��?.�EA�G.��>���.�>�G.��>�G�GWA�OZ�  TX;�u�X @P��X� @t3�ø ø �P�	�!X�3��؋l.�^w u��u.�^w u
�l+�=% r���
�u���bt��eu���
c:\drvspace.ini   Invalid setting in the DRVSPACE.INI file: $                                         ACTIVATEDRIVE �|FIRSTDRIVE �{LASTDRIVE �{MAXREMOVABLEDRIVES �{MAXFILEFRAGMENTS �{ENABLE386 |ROMSERVER �|CHECKSUM \|DOUBLEGUARD �|SWITCHES .|AUTOMOUNT �{USEMRCI1 l| �|��DA�y��Es���Ss��<t�N��z���<=u\��rW*DAs2����EA�<uEì<=u?��r�w>�� ����r*�G�w>�<t���Ϭ<=u�r�y����<=u�s��u@��멬<=t�� �~s�� =2 s�2 ='v�'��>��>끬<=t�� �Vr��\w�n��<=u�<t </u��<t�<F� t<N� u	^w���� �<=u��r�9B�0��<=u��r~= wy�t� ��>���<=ug�� rb= w]�t� �9B����<=uK�� rF�`w������= s8�����ǃլ<=u)� r$�E�<,u� r:Et�� = s�E�<t�	�ez�!��z��д�!��u��
��!����ô>�cz�!�DA*y�v EA������ՊD*DAr��:EAr�EA���硁��:EAr�EA�CA2���ì�� <Ar<Zw�<:uF���ì,0r)<
w%��ج,0r<
w���
 ���u�s����Ë�N��3�N�úUz� =�!s�Sz� =�!�czþ�z�2 r/<	t< t<;t<t�g �F���zt� ��� <u����z�Ëcz��z� �?�!Hu��z<t<
u��ð�Ëހ= t�G
�t:uF��G�%�G
�u�������<ar<zw, �  �~
t�H���"���.��> tS.��>�Ã.�su.��>�[.��>���=DStғ�u�+�� �˽ � ��.��dD�H�u��Mx�������u;�u������?������u����2�ă�@����������@���
���Mx��Ȫ���Đ�u����$Mxબ������u@�u������?�����u����2�ă�@�6%���ȭ�Ѓ������@��
����Mx��Ȫ����ƨu����$Mxߪ�������u@�u������?����� u����2�ă�@�%���ȭ�Ѓ������@���(
����Mx��Ȫ����ƨu����$Mxߪ�������u@� u������?�����@u����2�ă�@�:%���ȭ�Ѓ������@�w�	����Mx��Ȫ����ƨu����$Mxߪ������� u>�@u������?������u����2��@�x% ��ȭ�Ѓ������@���V	����Mx��Ȫ����ƨ u����$Mxߪ�������@uH��u������?������u% ��ȭ�Ѓ����	��@���% ��ȭ�Ѓ����	��@�q������Mx��Ȫ����ƨ@u����$Mxߪ������ꨀuJ��u����	��?����	���u% ��ȭ�Ѓ����
��@�[�% ��ȭ�Ѓ�?���
��@���p����Mx��Ȫ����ƨ�u��$Mx⪬������uF��u����
��?��B��u% ��ȭ�Ѓ������@���% ��ȭ�Ѓ������@�i���Mx��Ȫ������?t�t��x��֋�+�&�&�&��������� ��٨t$��������+�x�֋�+���������t ��������+�x�֋�+�����:��t.��������
+�xŋ֋�+���t�����������N�t.��������ă�+�x�֋�+���t��������0���g��Á�?t�t��x��֋�+�&�&�&����r�������٨t$��������+�x�֋�+����������t ��������+�x�֋�+��������t2��������ă�
+�x֋�+���t��������$��i�� t.��������ă�+�x�֋�+���t��������������?t�t��x��֋�+�&�&�&�����������٨t$��������+�x�֋�+����������t ��������+�x�֋�+�����X�� t2��������ă�
+�x֋�+���t������������@t.��������ă�+�x�֋�+���t��������8������?t�t��x��֋�+�&�&�&����z��%���٨t$��������+�x�֋�+�����&����� t$��������ă�+�x�֋�+��������@t2��������ă�
+�x��֋�+���t�������������t.��������ă�+�x�֋�+���t��������������?t�t��x��֋�+�&�&�&�������;���٨ t$��������+�x�֋�+���������@t$��������ă�+�x�֋�+����������t2��������ă�
+�x��֋�+���t�������������t.����	����ă�+�x�֋�+���t��������5��	����?t� t��x��֋�+�&�&�&������Q�
�4�٨@t&��������ă�+�x��֋�+�������� ��t$��������ă�+�x�֋�+�����w����t1����	����ă�
+�x��֋�+���t�������������t.����
����ă�+�x�֋�+���t����������
���Á�?t�@t��x��֋�+�&�&�&������e��H�٨�t&��������ă�+�x��֋�+�����K��4��t#����	����ă�+�x�֋�+���������t1����
����ă�
+�x��֋�+���t�������������t.��������ă�+�x�֋�+���t��������C���� �Á�?t ��t"��x��֋�+�&�&�&�����1��v��Y�����t'����	����ă�+�xދ֋�+��������C���t#����
����ă�+�x�֋�+�����l���t1��������ă�
+�x��֋�+���t����������� ��t,���������+�x�֋�+���t��������k�����Q��ـ������sZ% "��+�xJ�֋�+���t�������ZЀ�rF���ҷ ��.��dD���sN�����ҷ ��.��dDY�E���s
%? B�����s% � ��
두��sڴ ��낅�u
.�sut
��.�suu�����>�o�.p�p��t	���s�Ī+>�o�PSQVW���p�p  ��o�6�o��o�>�o��o�� ��o�����t�����6�o���>�o�ru ��_^Y[X���>rut3PSQ���6�o�o�&p���. p��r&�&�T���Tu��T� �� ˇۃ�r�&�&�T��T��o��o;th����];t[����];tN����];tA����];t4����];t'����];t����];t����];u�:Gu����ou/���ls�m�����������E�ֈu���T�����lPFI�D��ֆw���T�����l����+߁�?s�S�������ٌڎ�o��tNA+�S��S���r&�PIu��. p� �P��o�.p���>�o�.p�p����ې�^ ��
�yXz���s%ۋ�*���ƀ�6&����̀���À��"��ۋ�*���Ɗ̀�	&�����À��^ ��
�x���@s&������*���Ɗ̀�	f&�����À��W��@s)��@������*���Ɗ̀�7&�����À��(��@������*���Ɗ̀�&�����À��^ ���� w,��pۋ�,p��*����*�&��������À������?s)C���� ��*���Ɗ̀�&�����À�� ��s(C����@ ��*���Ɗ̀�&�����À��v��� s(C���󀀋�*���Ɗ̀�&�����À��H+ҋ�*���ƀ�&����̀����C�����*���Ɗ̀�&�����À��������*���Ɗ̀�&�����À��.p�p�>�o�&pY[��op;�orX��ru���QW����T��o&�&�E&�E&�E
��Iu�� p�T_Y� ��������*���<�.��> tS.��>�Ã.�su.��>�[.��>���=DStғ�u�+�� �˽ ��.��dD���u"��Mx�&�G�Ċ$F�u��Mx�&�G�Ċ$F�ڨu>�u����?�Ċ$F��u��2�Ċ$F��@�:���������@���h��Mx���&�G���$F�u,����$Mx�&�G�$F�ƨu����$Mx�&�G�$F���Шu@�u����?�Ċ$F��u��2�Ċ$F��@��ȋ��������@���
��Mx���&�G���$F�u,����$Mx�&�G�$F�ƨu����$Mx�&�G�$F���Шu@�u����?�Ċ$F�h� u��
2�Ċ$F��@���ȋ��������@�e�]
��Mx���&�G���$F�u,����$Mx�&�G�$F�ƨu����$Mx�&�G�$F���Шu@� u��
��?�Ċ$F���@u��	2�Ċ$F��@�U�ȋ��������@���	��Mx���&�G���$F�u,����$Mx�&�G�$F�ƨu����$Mx�&�G�$F���Ш u@�@u��	��?�Ċ$F���u��2�����@���ȋ��������@��Q	��Mx���&�G���$F� u,����$Mx�&�G�$F�ƨ u����$Mx�&�G�$F���Ш@uC��u����?�Ċ$F�x��u�ȋ����	2��@��ȋ����	����@�f����Mx���&�G���$F�@u,����$Mx�&�G�$F�ƨ@u����$Mx�&�G�$F���Ш�uD��u����?�Ċ$F����u�ȋ����
2��@�[�ȋ����
����@���>��Mx���&�G��$F��u&��$Mx�&�G�Ċ$F��u��$Mx�&�G�Ċ$F����uC��u����?����C��u�ȋ����2��@��ȋ��������@�$���Mx���&�G���������?t�t��xً֋�+�&�&�&����/��� �f�٨t������+�x�֋�+��&������Y�t������+�x�֋�+��&�������t+������
+�xˋ֋�+��t���&���&�������
�t-�����Ċ$F��+�x�֋�+��t���&���&�������#�Ł�?t�t��x��֋�+�&�&�&����������٨t������+�x�֋�+��&��������t������+�x�֋�+��&������t0�����Ċ$F��
+�xƋ֋�+��t���&���&����d��1� t-��
���Ċ$F��+�x�֋�+��t���&���&����/���J�Ł�?t�t��x��֋�+�&�&�&����������٨t������+�x�֋�+��&����p���t������+�x�֋�+��&����_�� t0��
���Ċ$F��
+�xƋ֋�+��t���&���&������X�@t-��	���Ċ$F��+�x�֋�+��t���&���&��������q�Ł�?t�t��x��֋�+�&�&�&����;�������٨t������+�x�֋�+��&���� ���� t!��
���Ċ$F��+�x�֋�+��&�������@t0��	���Ċ$F��
+�x��֋�+��t���&���&������z��t-�����Ċ$F��+�x�֋�+��t���&���&��������Ł�?t�t��x��֋�+�&�&�&����������٨ t��
����+�x�֋�+��&���������@t!��	���Ċ$F��+�x�֋�+��&����y���t0�����Ċ$F��
+�x��֋�+��t���&���&����T����t-�����Ċ$F��+�x�֋�+��t���&���&����+��	��ā�?t� t��x��֋�+�&�&�&������@�
�#�٨@t$��	���Ċ$F��+�xߋ֋�+��&����D����t!�����Ċ$F��+�x�֋�+��&�������t0�����Ċ$F��
+�x��֋�+��t���&���&���������t-�����Ċ$F��+�x�֋�+��t���&���&�������
���ā�?t�@t��x��֋�+�&�&�&����1��[��>�٨�t$�����Ċ$F��+�xߋ֋�+��&�������,��t!�����Ċ$F��+�x�֋�+��&�������t0�����Ċ$F��
+�x��֋�+��t���&���&���������t-�����Ċ$F��+�x�֋�+��t���&���&����r���� �ā�?t"��t#��x��֋�+�&�&�&���Ċ$F���p��S����t$�����Ċ$F��+�xދ֋�+��&����r��@��t!�����Ċ$F��+�x�֋�+��&����U���t0�����Ċ$F��
+�x��֋�+��t���&���&����2��� ��t-���������+�x�֋�+��t���&���&���������Q��ـ������s\% "��+�xM�֋�+��t���&���&���ZЀ�rF��������.��dD��sN����������.��dDY�C��s
%? B�����s% � ��
���sܴ ��끅�u
.�sut
�,�.�suu���� �>�o�.p�p��t	���s�Ī+>�o�PSQVW���p�p  ��o�6�o��o�>�o��o�� ��o����t�����6�o���>�o�ru ��_^Y[X���>rut3PSQ���6�o�o�&p���. p��r&�&�T���Tu��T� �� ˇۃ�r�&�&�T��T��o��o;th����];t[����];tN����];tA����];t4����];t'����];t����];t����];u�:Gu����ou/���ls�m�����������E�ֈu���T�����lPFI�D��ֆw���T�����l����+߁�?s�S���������&�tNA+�S��S���r&�PIu��. p� �P��o�.p���>�o�.p�p����ۋ^ ��
�yXz���s%ۋ�*���ƀ�6&����̀���À��"��ۋ�*���Ɗ̀�	&�����À��^ ��
�x���@s&������*���Ɗ̀�	f&�����À��W��@s)��@������*���Ɗ̀�7&�����À��(��@������*���Ɗ̀�&�����À��^ ���� w,��pۋ�,p��*����*�&��������À������?s)C���� ��*���Ɗ̀�&�����À�� ��s(C����@ ��*���Ɗ̀�&�����À��v��� s(C���󀀋�*���Ɗ̀�&�����À��H+ҋ�*���ƀ�&����̀����C�����*���Ɗ̀�&�����À��������*���Ɗ̀�&�����À��.p�p�>�o�&pY[��op;�orX��ru���QW����T��o&�&�E&�E&�E
��Iu�� p�T_Y�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     SRVWU�Ȏ؀>�� uN� � �Ӏ�@*DAr:EAr2SQ�D�!Y[r'
�u#SQ�D�!Y[r
�t2䓲���ҋ�
�uƇC��� 3ۊ���
�t,A2�Ƈ��C��3�3һ ��������Ku�3�5�7�9]_^Z[�SQRVWU.�>��r�� .��>��"���؋�3�&����u�� ��.;�>t�H.;�>t�&�G�Āu���t�� t�.��>&�G��X &�G
��^ &�G��` &�G��b &�G��d .��������.���.����.����� ��\ ǅZ � .��>A�>�v >�V�D �>�F >�N�ى�D ��F ����R � .��҇�.�����A.��҃�s���,�]_^ZY[�PQV����3���9��u9��t����^YX�QSVWRU�ߋ����2Ұ��[Cu&9ou&9Ou&�w&�:�s������]Z_^[Y�QRVW��3�� ��u�?�	.���>�t^��.;DuV.;DuP&�G.;D
uF&�G.;Du<.�\>�F.�D
.�\>�F.�D��?t����.DA,A��.���A���u:�s�Ѓ�⊊�_^ZY�                                                                                                                C:\DRVSPACE.000  
.�����o����3����# &�� .�J.��>&�� .�L�7 &�� .�N.��>&�� .�P�( &�� .�.��>&�� .��PQVWRS���#[Z_^YX�2���{Չ}�P�`K��?��D��>  X���վ���Ԋ<�u�AS�xՀ| t�\�x�,A��2�ۊ��A[$A��ՊD*DAs�D*y�r�z�2��6EA�Ģ�ՊD2��6�Հ�0�&�՘�6��00���QV��մ�}Վ{�3����s	���>�>WQPV�)��> t7<u^XY_WQPV���BL�)<u��> u�^XY_WQPV�q)�����RV�G�<	u�?^Y�D	���W<t
�u.PS�����2��h[[X�	t�<t�G�P������X^Y�D<t
�u���| u���DA���I��DriveSpace found a problem on compressed drive @.
To correct the problem, type SCANDISK @: at the command prompt.

The startup process will continue after 30 seconds.
To continue now, press ENTER.
$
Drive @ is too fragmented to mount using the current settings in
your DRVSPACE.INI file. DriveSpace will adjust these settings,
restart your computer, and try mounting drive @ again.

To continue without mounting drive @, press ESC now.

$Compressed drive @ was not mounted.

The files on drive @ are currently inaccessible.
$
DriveSpace could not mount drive @ due to problems with the drive
or with your system configuration. You may be able to correct this
problem by typing SCANDISK X:\DRVSPACE.nnn at the command prompt.  For
more information, see the README.TXT file. (There is a copy of
README.TXT on Setup Disk 1.)

The startup process will continue after 30 seconds.
To continue now, press ENTER.
$
DriveSpace could not mount drive @ (X:\DRVSPACE.nnn) because it is old.
The startup process will continue after 30 seconds.
To continue now, press ENTER.
$Drive @ is only partially converted to DriveSpace format.
To continue, press ENTER.
$DoubleSpace drive @ was mounted read-only.
To be able to write to drive @, you must first convert
it to DriveSpace format.  For more information, see
the README.TXT file.

To continue, press ENTER.
$DriveSpace could not mount drive @ because
it could not find a valid DBLSPACE.BIN or DRVSPACE.MR1 file.
To continue, press ENTER.
$
Compressed drive @ is currently too fragmented to mount. For more
information, see the README.TXT file. (A copy of README.TXT is located
on Setup Disk 1.)

$DriveSpace could not modify your DRVSPACE.INI file.

$DriveSpace has adjusted the settings in your DRVSPACE.INI file,
and will now restart your computer.  If your computer does not restart,
then restart it yourself by turning the power switch off and then on
again.$PQVWS<u�Q��
�u�� u������u�-�� �� [_^YXÊC��$t��@u�xմ�!���SR�@ ��&�l ����!
�u&�l +�;�r�2�Z[�QV��A��!�O6��!^Yø����.�>˹����3�3�����1���ر���ȃ�&��>&��>&��>&��>.��>&�>�&�Z ��N .�>w> t�� �����=Ju
���t���tO�c4�u�Y.�>w> t��%���h��.r�.+�>.�>v� u.�>.�> A uS��u��vB����8�+�[���.��>�) �.�>w> t�����.�r�.�> A u�):�vB��.��>�.+�>������Y.�>w> t�����������+��ǋ���+�������.�> A t� ��u�vB.�r�.+�>���+Ƌ�����s���u-vB&)?&)?&)�>&)�>&)~>&)�>&)�>&)|>&)�>&)�A&)�A&�?&�4&��>  3۹ &���> t&)��>&��WA t&)�WACC���!.��>��9F u�>D 2 u
�F �D �B��.�>v� tP�.��>X.�>t��C �.��>��7 .��>&� � �VQ�Z�p>+΃��.��>� �&Z��&M�5BY^�P��@t�Ǳ���ȃ���W.�6�>.��>���������_&��>��&��>PRVWU&��>��������&+�>�&��>&�>�[]_^ZX�+�&?&b?&�d?3۹ &���>�t&&E\&�U^CC��ÿ��3ێøJ�/��@uJGtGO.��>���;�w:P� C�/<�u0�C�/.��>.��>XP�ظJ�/�tX;�u��@t
.�>t�.�v��.��>&��>� �! �& �+ � �0 �: .�>w> t�� .�> A tA&�xu&�|u&��u&��uP�ȃ>5  t95 u�5 &9`Bu&�`B&9�Bu&��BX�X�.��.�	���R�!&�>	�t�� ����     ���������            ��Uuk
�tg�.��.�EA2�*�s��.��.��+�.���.��  .��.��.��.�DA,A.�!�.EA.�#��!.��. DA� �~ �� �?�o�.��>&�.�#�&:v>.��>&;Gu.��&:Gv
.��& G�&(G&�.*!�.:�s.��& &�_�.��.�EA&(&�_���.��>&��ˌ�&�_�.������2�&�:�r�Ћˌ�&�_���u�.�>��u�����&�G�D&�G�DS&���&8w�ˌ�&�_���u�[��ߋD&�G�D&�G�\�D.��� 넹 ��A.�6�$.*!�.:�s7����.�!�.����.���A.���A����2�.���A�����.�>� t*.��. z�Q.�EA2�I��>.��>�G������Y���.��>&�_�X.�&!��.��.;�tV.�X ����- ��.�����Q����P�P�P�P���E�E�E�Y�����!�A&�����X��ðX�&����QC�W &�&� &�C��Y���    c:\drvspace.ini 
MaxFileFragments=����>+��>='v�������2 ��滵�����Z ���<u�������Z �����A$a���C3ɺ���!r8�=�!r1�����
��梙溘� � ?�!r;�u�>��u�B������!s�{��r�랺�� �>��
t����� @�!rޡ���5 ��� � @�!r˴>�!rŸC� ����!r���!����&��Z �8�� 
 3��6��R�t���X0��溙� @� �!�.��վ����D<tv�<�tp.�xՀ| t�\.�x�,A��2��.���A$A.��ՊD2�.�6�Հ�0.�&�՘.�6��00.���VQ�ڿ�ڀ|u��ۿ�۾�չ ���z����Y^��It�z�� �5�!���t�@ ��� �SO����@ ���r 4�  ��PSQRVW3��ǿ� &�E&t^�J�RM�IC�/��CIuM��MRuG�>�@��@&�E%� =� &�Eu�A� ��A%� =� u�%` =` u��>&;Ew	�_^ZY[X����      V&��> t&��>&�6�>�3��޸J�QS�/^�&��> u���&��>&�>�>�� ����m'�&�C-mmmmm
mm�U*�߃��� ��C9t���
���u�/��&��>�h��&��>&�>�>�� ����������E'+ǉ}'��&��C))E)E)E)E)E
)E)E�U*�߃��� ��C9t���
���u��?��ǉ�*&��>������> u��> u�,��+r��A.�NB.�>B� =�NB�!s��ظ ?� ��>.��>�!s�� � ��SQ�CJЁ�P�;�Xu���� >�!� =�>B�!s� ��>�ظ B3ɺ @�!� ?��.��>�!s� S.��>��C�?� t���[�}��u� �u��u� B3ɋ�[.+�>���?���!� ?��.��>�� �!rA� B3ɋׁ� ,�!� ?� .��>�!r%� >�!�r�.��>.� A.��>&�H �� >�!.�&�>���SQRVW����>&�D 2 &�F &�5 ��B�`wt3��ǿh &�E&u�� ���RM�IC���CIu��MRu�&�} tw"� &�E���� ;�u&�} tb�ȋ���#�u�� &�} �w��� #�;�u&�} tT�� � A&�M
&�U��B��B&�]&�M��>&�H &�J &9L t&�L �/&�=MSu�&�}FTu�&�} s�&�E�����&�E� �&�E
��&�E�u���>�< � ��3����� ��- ��>&�&�U���u�bB�ʣ^B�`B��>&�0 �����t���� ��_^ZY[���� � L�!                                                                                                                                                                                                                                                                                                                               LE             �                        �   �       L       �      �               �                 �      �       �     � 2                                                   ;  -      E             �                         DSVXD    �           �    �       O   �  G  �� �' � 1 �W ' 2 o ' ! t '  � t' $� m h ( , �, � � �  �  �    _   h (                                                    ��u��  ��u�u  ��u���3��  �t3��.  �  �t	f� @�  3ɇ  ��=  ����M�w��wr�E;(  sf�  �  ��f� @t��3��r�S�%$     � ;  ;$t(�   u��   u�s�f�fC��f	NC���   ��[f�e,��f�M,�P�E�=  ���Gr��	�r�G�Gt�G�u�,  �   �wXÇG�t����   ��s�=  �3�3҇W�t�   f� @3҇�t�   3��G����   ��R�%$  Z   �f�`C��f	HC��ù   �   f�S�������  �   �,  �0 ��  �   ���    � J� �        ;    DSVXD      �    W                                                       X                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           j j� �  ����n   �  ��lW�|$� �  _� �  �sf�F R�!   � �  �~8���N��G��������   �G!�(  � �  V�t$� �  ^��l��� �  ������Љ  ��  �   r��  �R������Љ  ��"Win386 DSVXD Device  (Version 1.0)  	DSVXD_DDB                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                � J�#;�si��-D�%������ ��~��ر����S3�S�PKLITE Copr. 1992 PKWARE Inc. All Rights ReservedNot enough memory$� 	�a�!� ����OO����������FF� ��� �2�����;����<����A����c����d����e����f���r���Jt�s�3�3���Jt�����Jt��Ӆ�t��Jt��Ӏ�r��Ju�����.����
t:3ۃ�t&��Jt�r��Jt�����Jt�����Jt��Ӏ�s.��,���V��+��^눬Ȁ� <�u��3��Ju����Ӏ�r���Ju����Ӏ�r���Ju����Ӂ�� ���3�� S�؋ȋЋ����� 
      	          	
� � - SYSUt �ility � � ���, ����  ��،��|�&�� ����!�*rT�>� *C�P�7��`4r<)P +r6� �=r+
��&��r8P @	r�
r�0 r�
� C�!� �	P�MXP�_X
=u3�� 
P�L�����JA/��3���*5�/ �#C3�#r�A� ;�t������   t�= �� 2��\Q ����\YA��G�a�3DA7U:TuO�) �&, ��rA
�W���6&  6��sY_�)� G� &�*t�� �< u�FG��Y^e��_����T��,�=\uR� H��� ��Nvs�>'((- t��Ų  =�~s���?��@�N�`
�n;�t� ���>
u
&(P2C���P�<[I�%X:�Lr6�ȴ@K�)�J D�uyE�Lu�?Wb�p�!���>�3
�
��X�_T�s��g� ( u���W� ��� �u����B�_��s$�)@p0)��=tAF��r@�� ��  r� �<�>��(P =  ��� �w U��u#WV  �6�����3��\ ^� _�� ���P�� �"�&�J�5 ����2�SX��Su�a E�B��u�(���Zl
 vP
�ì��À�C( v���
�u��� �&�}�\t&�E�\��#)�6 �3���'Š�����{@�* &Ío.״'�è	� �>��u �,� �@���� ��_=/�At@��� � (�# r �sr�%P�\�����J@:XH�Yx�)PD�`;��`;�����	%�u�� 
U�6 �,���t�>� �ԑ,N)J��?>��c'T��@Y��B~u���B�'�B!�R�G��UO>O�}[�S�
n���qI�oÀ�<�t����@����P��r
�À@t��$��J3�P@�/����MD�A(r��

I�ÊL�ŤD�=��S�4��r#EQ!:t@}����-��8%2���I	Ir�m�� 	//
����!�� �rM��2EB��D s� s��`I��Z �	1� �`$d�>�c$u�B	��ь� �*���� rF��R�5�Jv6r0�1< t-G�>/�I2�>dʞtDfs s�U���V��r- ��������;�o��Ы���T
��Ѱ) �
�Xu���s�^Ë�� ��r��s���xr�XmWa�t�
����� �r$�D�E��&����-���M�U�ġP�V�
�$3��<,r�+@ȋ��}9P`Ms��uP�����?Q.��*)h�].= �;�s
�̓�<�L=��S_[�
�.b]G�  (U�]
���uPR�H=�U�E6�ZX�r�@�Wu+�,�vH��԰|)�� r��)������"�>T���� R���i���<�t�uv�6  ��>�� ���u�p"�|� u�`��RJ�
&�'u��'6u4��x,F�OG� ���n6z�]������N
� Tl����RZ�ڎ�r!  {P���`P@��D���P���ý*���� ��u����E�i�@$�u!�P! ����|����,� r0"�r	�r�����R� �~�Uu}rzhUx�:z�� rf�� {(0�{t#�^ut(�uvt�t���N`�!����P�����,�"(��-����@"�6��ᣖ���
d���s *�db�e!���W
�UR��#MK��u"�$���4 ��46�' �>FT�H;4�P��P �����@��8 r  5���G ����� r"��"EU�ZbUUowUQYYu�(@H���
 ��)�j%H"����/� ��r �0����7J$"t��!� �
�<!�y.r,�6�,  ��"<���O��!"��l�!y�� �@s��	K�gI �P�<��U��!M�W�gt��䵇�������2ĺ%�cV�D"�i" ��V��<u���s,��0��J h�6��>�ɤ$�n!E X�Rra ,0�� ^6�u����2��I���%�(3�L%% �<J%!Jl���ls />�u% (�á2�  ��jH H3��q�ȡ7�&1�
/4�+�3�9.��("=�w�6��`��-�D�*� ,!P�������2��΀� �w��u� ,�.��eh 0A*�#w�/ �� QD�((iuA �u�2��s
裄������SY�v[iê�Z�2�(@�&��$�����G&��3��G�������F�R�� &��� ��r&��@�&�������H��$	��85�&�U��$)P�&��K&YJ��M�'1�aV�P!U uI*�\4E1R�@&�
�ngTuÍ��>��6X�=�ȑ�J 	���Ƌ�>T�2N rK�+�_ �;�Kt���zPC�R"�BjI �K���D �E�Ku
�|7u� �2H �j(��	Ar�;�r� ����r�)�[���b�w'P�Y s� �r��v�����VU �l����%B��Kp�
��%����x�%� 
�&X]^â�����*���t@��@�`T�t\�?��|�
��
�5E�-�%�!�o(0Z<�u�
�]r���
�dU��%��s�R@.B��QWRS�^�櫰��U
��r���o[ZY_�_2)G�E�6U0��t)��<�D	�HE��H;q�3����>f�NxH�7�@�r;>	u	�6b	$F!;6���v���}P��o�j/J) �h3�3UU]	�L��PIU��E�K���Mā_X
����	)
�6�
 $i�^�g�ێÐ\Ό��؄s	5l�"\�`��5u��~w�L������6W$����H���E �����r%�B�8�>ppt
���`
�G�  ��%������Z�K���HH����n@� Ä�$  �#�$�.��D ����r��Tv*tj��H�w��F��;�Q�{�%(��T`�)QD��5�G�7@����=Y;�vA��闊I+H� 8��Va"_"w��fMV;�sS�34�4Vs*a?YY��'C:�E�l��H����gu!P�P��>8IC���@;��X�t��I&n����b�����!sB��43� �n�(� ���� �؀?�u�@`��G���M%%
.
��txp�*�M�yO�n�{�X��ؿ��ڹ�rE�%.*r8��8- t)�B���g	E��Z�"��r|�Lw�PA�Q�y���y* �����U�3
@�y�[r=��R�y j�tE[���	�X�&3��?KH0�
0@�� ��M����� Es��u=���������s�3�*����&v�������!�+��f�shFQG`�6C��i{+	8�<02	H�8uHe�~�����d's�eoj�  ���R�!3�&�O!&�_! ċ>h�  &�GC @t�u �&8u
&9GIu&�I��X��ápPP�� c�	���/��f�}<AdUtNh@H@tC�K}�!�E��r#�	�@G:�4��2!��s��`0 ��v��*Tr.-��Jl~8v�����zx�f���b�rR�6�Z4��\D^�8 �]�Z �.��^� ���aQ�>j�x8�w�� E��� V�h r	�� (�9��^����bV�ƕ'l���8�XV9�a��������!����+�<s���� �< ���<^�S�
;6jr�w]+��N�tH���``#t+�Q9P��P"+�;$sWD7.I;���/� >��3ɊȊ�2�P��@�R��s��2W���ѡӆģ�%������ts7���[� ��
�t:  �t���V�ذ\&:E�t@����&�����
��u�� V�Zp��<I
WU7.hIl �C �O .:��	~�<t	)
.O��l.�!t (��o��O� �.�C �O��.��Vi.COMJEXE W������WPo-O� ��4"G�F�ǧuE!����obR��l_Í6e
���*
�	;�3�&�E, ����VQ�Z^tO2���&�#hy�u���;P*   F��  Invalid dr  ive specificatio nExtendeErr or %1�@@��@�D  
	 D	 7LP  @Too many parame�=rsRequirD� #issing~UPf^P�8t noc�t.ctsey��yu��y, ( -^ .z /��   � MCopies MS-DOE)S�ysYmY��il���Xmmyl�qprwt�a
���k youP��y.
e^[1:
][�th]�t#2: ? �S;o��lo�=D of�y�bF N ��@��e
�r)S�bc�d&.GIn�E0 �2rs� t/�0 ��+0
 (�M�  r 
 �  �  �   � <  (F(NbroomxS���d�s��nϠ<.`(�U6�#-So
��Bund)dtransfe��g^fau΢lt�C�*A�NU"W9)e_ajuM,��etousaU�b#&B��adfrT��s�rc'$��c+o�Lm�E��+targeo/�EC0ld�p��MANC2D�/�.�1P�I�ufPAie mzo�ry�-��� �   0  � j  ��&  � �%1���nTw=kW�� Y�tw�еin��'1{' !�!#N["g�H�j�]V:$'�SUBST j�ASSIGN^ed�1SE�ixV6�Ub�s��� ����  C  !Pres��y key�c(eQ�u4.� 5���0�P  SRW3Ɏ�3��.�v�3��>iJ۔(�)&AI
�=�J*$")m�-S-0.�M�F�$12R�T�
 ��28)�(�6%�%�:S>R *= �r_ %Z[X���
��V. Fc�!r$ĉ6F~H^X@d�D�/1"����&1�n��
PSQUW���@��J�6Oj��@t#�u!.��"�rZ�x
�2���{�*
Z�u]Ye2[� �N�HV&2>,>w�� s�Y�l2��8t��� r;��i� �u�&�-��$e� sU�j��Hڑ�	 �����WPS���eٰ��+�K��[X_-e�-OAܦ��Z(OUP�\&�XX���B�P�u����� D��UQ����Y�R�ةȘ
�;��"]q�'� � ������ƀu��M� � �OW�>F� &��t&:Dr'w��GG�� � LP3ۓ��6T� 
��	v��7�0R cA�u�t9 ��|
,u�6]AJW�"�� ���3��T���e �!�%�� &8%8e` t:�uS�
 s�BIu�V���t3M�>�u+�DfA0���<0* ��64��>O(�uB4IOO��  ��W+��
�_Ys�e�Q
R�ʊ tu%#�^��R�	U�:�ɂ�<pQ
m�DS�|
��[n �{ 4  rY_]^���*pH.�0�K١ P6��X��VC��@P`j���q�
��C���VS3�Uw����2�@��%��tu��È�=�='�T w"!����7)%/�p�𽄪>��� �T ����(r㼟�+��u)RUQW ��/<�Xu	����*_�\.�� ]Z�o[^�	x2����I�"�\G�c'�t �P������ �t&�M�	.85uE.��d-��}&;TR�.�	II��������}�2� 0FG�L ��3ۀ �u�; ��-CC�CVPn]3҈ %�D	:�v*���4��t
 %}| ��u�E8Ls*�*-ъ�$HS���A�AaB;�u�Uu
��Y#Y�,B�j�K�(��u��U�Q_Qoˬ�>��9�s�rq�D��]60u	xPA�Y�s�EPd���@GA��+�DR����v��$����x��P:
�t��*;Q�b ��� r[+Zd��[]|< >+=;" .�K%��2.�>%@�NSD*��%1�%6���%;�%!@�6s�	S&�&:
�\�#N6M@%SWU�UU�L%   uC���r<�*t7�[n`u���& AtN�.�<=u.�C�b�	��C�NWB(HP���Q%t��6`�</t6"hVGu�T&�G�.9�s.���C�C�2� �icu�`��(@� ��2�CS�('��sA4����,,4U�,
	@�6]66 ]P_[.�Y�5Q	��D�b�F%��P2�(��.��E����u	D=�P��0�� X�X���UQl �s�o	�Is P� ����.�.S��WY]�&�~���E��E�GB)��rJ&
��P�O%+�.M%Xt*�Oz&�
|�:|	|&1 ��&��Nu�"�q� &��m
����W�}>Pd�&�ec��&�X<��g�U0yM�Z<u���P<t���<�><T�u7�@8�T/�]/+
�
��9P&�G�G�g�	t�j
�{]y���H�% � S0��yW��̦�K�_H�%@�A��.v���.H�.�>+u&��\�
/ t
�ї �k��� uEBiX~.�(?<:u�P:��7�sFF��H��VR�� �(��r-Q�.���Z  ^�<�s<ar<<zw8$�  �4SW�>�%.8tPQ �R�e�»��� �r�!ZY�]��E CC,�&�_[E0r��<9w,0��,���u���	(>�&0	URV��<a	�v�MBt�S�q�ti��
hu\�A��FI�	�RFE$&�EFKE*�9@t1� �A�A%"a�TO	O�\`U:o0)�I��^Z]�WV� �>M%g��_)$�8^h_�?z�2��)X��
�-��\(`sGF��.�F%
�2G�B%^_XA	PP �'�qSQ��%�1�	�	�C��AY[�R�N8�r,.�|r:����� � H�,`��O�P����*Z!)Y��"��S,�qt��	N�	pN��<tq-�)<
t% �&�}r3�&�]��a9Y�	C&:R�!�/(�6�K( ��<[ �6<	t2<,t1u��� F:��eR�CM
[S� KʅK K �T� � 7�.U%;�It
</�ya
*� @�VSI'PQ�URWU3���P����]_ZYX���G]�Ia)
��
�t: �r:Dw\�+��[^�N� A:�\IO.Mb]
MSx!�IBMB�|λ��6; s;]6J � :P?]�Cx.�	:RCDRV GSPACE.BIN�;�.��H���[��Ƣ	/?vNO NAt ME  FAT12��	6���� �{g	$
��$6MS�V�B �(C), %yright P 1981-94 Micr��osofrp L�eKd�� c,al - Prb�"ty��� /Alb�MslQ:}v5c�dή �+pl@2Dq,�ŵ OIOԉ+/ ?�c  ��<�b�5.0 �9Q���
$� �)n e�3��м |�x 6  �7VS�>|� �� ��E��|�M������rTy59|t � |�|�&|��||G��PR|�IK|�  $|�
( �H��	R� � �'�(.� r��$ �����}�u
�Y  
t��}B�^�@�D�X�� �HH�|2��U��ZZ�YVPRQJ"�:Q�XT YH� �	 ���.|�$K��4�3�  p: �)�� �����;�s�6 ��O|3�|R�
%�M|Hn��
�P0��
6�ʆ�) Q�6!��
Non�-S]�6�e��Repl1�a�Y��pa��when�hl� l,���лU� ����@( ��Cc�^�d��PATH=Ax,SPEC=' �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        MZ�   H���    ��R   PKLITE Copr. 1990-92 PKWARE Inc. All Rights Reserved   �     ����    �                  ����  ; r�	��!� Not enough memory$-  ��- ���P�� 3�W�D��ː���S��- ڌ͋���������NN��+�+؎Ŏ������ 3���� �+����5����6����;����]����^����_���r���Jt�s�3�3���Jt�����Jt��Ӆ�t��Jt��Ӏ�r��Ju�����.��a��
tu3ۃ�t*��Jt�r#��Jt�����Jt�����Ju����Ӏ�s.��q���V��+��^���Ju����Ӏ�r���Ju����Ӏ�r���Ju����Ӂ�� ��뼬Ȁ� <�u�[���3�����Î����&����Ò���ҋ����S�P�Ŏ�3��؋ȋЋ����� 
      	          	
    :  �Y����м �`U��V �T �P ���R ����  ����،�+شJ�! P�X &�� 2� 
�, 6�Z �R� HF�< u���V�	 @���^+ދ�J�C���I+��N��� ���6� G6�>l � �N�6�FG�T��3�	)�
�+�P�o �L|9�U��� U |��v�� 8A��]��F��9��~��1�P�	.���� ��6X.��]<| �l���e�c�
��!`�e X`� � (�.�F�S�
��*��	�
�Pz��P�<���*8��t,�8+�$���,T�d�CI*c��X(��tQ�4d*Ci3
j
U̸X]1?�K�0u3���2R�> e�t� ��P��'Q1'J�!'u�l
ŋj/=
t
I=-=<=�,����L	!P$�;I��9��6��Ņ	5�� E2�,#�H���>(��@�C��F�B�
�D"( ""��Uo��RW�8��9�)) � �},V� ~!u7�^��W 
��V�����v����M��^�?$�*��v�@7��/�<��9HPr�� +��Զ\��/�^�  ��+���+)�+@ ���@�P��� H�o��0��@Zk�@uk�& `�ӎI�4AI�/E�u�E	E�E僰&/=B��@+V�d"��U��؃�R�v������K
@�.� �,C�*V�F�!@ }�*��B�E���~Q��r�.�$(�F���-�D�@(�F@�/����%f������j9 u#�n�?+u��6kF���g�bhnGr�-,v,s��$�,�y9,|,�)9,}$�,u^�,�,NJ�,�$�N�,�,�i�,9�C�K���%���-K�K���C�K��nK�,�,)��$�,���,�,	�r,�$�,��,	nJ,
,	$�N�,�,�
m�,[�,:�	M���* i,�P(w�v�����AP
�~�4�������~� u����D����	�_�l�~�8 �!Cf�,�>k(�:ul"%��""� ˠ�F�{�i����0���yF����B�tٶ����t �n�����N����r��w-RJ�'�)�!��R��J)�	��� �髰�7f�t;�4eb\-t&���t��tt
)M��!��y�D�F��
��^�?��� ��F�<+t<-u<n�b��� �R��
�	J5�����G(���
"W�uYhԧ���BG�&V��;����l}ll�,�:t:�)� �+��aA�j��G' �@��^�)�OB�@
��Q��Ӄ@@Pl��l>\jGD0 �!��,@��Q};+����nu<sJ�ie"M6H�	pul�)h�7'�Z	�+)��p��N�H�N��@t鋔v����p`��	� ���v��HRd�Ɩ��+���jb���-�"�1�8S�4p��(*8�K,B-��^���21Vt?t�b*u�_�����$ 	���'�~^�ܗH� ��GG�{�6�6��)� �P��?5�?? 7�7���$���N�*��S^@���)�8]H�&��b�2���e������r⸕����
��ԏų$^6���Ott�o�t�A��tIt��et��mt.t�t�l�*�#iC�(.��A����S�DKDl�>� �'�N���F�\L�;\
�Y�Ӎ"Y��A]Y�F�@ � �LG �׫"�:��G��YX�nTP/�"
r�\gs#e�b�'bN���6k�H6Xt4p u��6"  ���% ��PQ�� L����f�*��F��J#!!��HE'"0��K\�!��\�0 Q�L�Q>G��W?��G?�]JGG�!V�1Kx����	�t2�"E�>b�BB� �&%���@t,
u%Q	�}W� �V� �� 3��33
3�3� �$��)"8
5�*�����B F��
�v��BP� ��~�s�H�슇/�5P���t���H:&��5 3'r��(�����F���m�����J���	�|��h�ES�� ���
 �L <<��<u@,�%�P=��u���!T��*r���)l����"�y����uFWS#W�> ���%�t�R8z ����6��z�����ELuRNL�$?�����G�GܼG�G��Po��� �AoF�"�m#�FZ�"BT�Q��tv`��7�~��G� ���ǆz� ƆZ� ��Ͷ.���F*�����#��Z`s�d��YPO��|�zZ�M�� ���.tF�$t?��HV9�^/X@X���!�N�`��������u1F6B��6�! ��eZ��8�q�
u�uV� ��.�yp!�3��&�>� 	���> g�'�O��t��r��t�����X��Ga���[�/'�TU�|�nH[eJ��S7�F�	����
�����$"9i$$5��0"!��	�r�Hu�~�&� �k-�#�%�l0���6�:�G�_%���� 	$�!z ��W7��٬4T����g \ 8?� ��Vǆxb��@R�B� ���p"� r��.��B�Ğ&�? Z��&8w��Gr�:D9G:�0�9���H1�^�`�K� ��|�����D��t��&F8B���}������e�Xj�~�����e�F�n���F!��Q%� D%�����y����F���T��	D��@���^�&�W�$巉���G� ,H��ԗg�(K�Vz�sL���+��D��CL����D��6�0�k�)
[�#���hC��E����`s�ht�U��) ��UEu��v�Y��o��u0��c	�rP 9QRSTUVWw1[��0��_^��][[ZYXϐ�S  ���FH˶[L�B]||>+ =;\WV���A��Hu�<^V�  3ۀ<"u��
�u/�=�@=�=t
=	)(	u� �F��VQFB%�Y^N�I;I 
FI�^
�u�_��2( s�S&�&:s	 �[��6USWU �]�T u>�� br7�&t2�W8�����"	@AtN��<=QP�C�\ɬC��NPJHU�Yj���6W�/t1L �t>uP&�G2��9Fs���CC
�-� �fq2^�%@�2튩��CS&�(f�s?3��+,��3+*]
	@5Tz�5
5 ]_[������ ��L�N��PBH�� u&�F��1�u5� �P����� X��KX�	P��5 r�& P
�P�W+�UX& WW@t	�#���f��Dí�B�BlUQb��O��oPP)�sL ��P�-�.[�Y]�&�~ pؐE��E��m���rBm�3mu#�|�:�zK�!ݮ&��E)�g� �c��
��W ���>L&�e* [~&�EX<jQ$	U M�Y<u�O R<t�<t�<�%=<u��@�R7.�].+6�
u
P&�Gt�2&	t��5�x�� � _�� с}�PSRW�
ġ��` ��_Z[X�� .�Q�i�>��!u��c��s*M?�@� 8�s���#�� $V�* t	����>�M� 6 ��X�PV�
�t@@<:u�|f��c �sFF��^#VR��%�r*�0 ���Z^�<�  s<arB<zw>$��:S 
W�>��t	8tu�e��»���}�͡ !f�]�EC�C,�&�_[�4���bo�	�	�F賀�GV3�3�S �B�r92��� ������ r,�ڋ��[��	�
	����	RՃ� �r���[� [� t
���҃�&�bwc؈���� F� t^F,�u&;L��r6&;T.�w(�w ��1||	
| ���	��u�L�{ `�; H`$�4�	��@�lӦFCuAt��11�1t`1
���^F6 Ü�u�Ýp�� ���<0r<9w,0�!�	��
�uDJ<"Oa>Gvӫ�

G H�-�0 s��}S��q�
ʿe���Ȇۅ�`��gURV� `'pr:���"L�tahXn�AtkK
uZF�Z&b:F?�6�PFE#CeKFHE
9 �7@t&�G  t�
P"e� �	��M����:t�p�S�^Z](:SV� ^��� ����$��(
�M�Le��Y�"�R�@���t,�uB�ȡ%	9�� �#u���U� �R#<	 #��ds��l[^ 2�S���H�J�Pȍ6e<�t  RP� 8���!XZ�"ÿ3��;�M�>��* r�t0<.t,��<-t&�"  ���r� ��
 ��  �u�r�F뿊���F���pTV�U�
�C�*�� #D ��F�� ����6Y��	^[�� IO�$t!� :���FCC�����ts5A�����J%@�2Wm>'0m��W u ��.^_�9>��-e�%X*C��
sYGF��&
�N�G�>�^_�HX	P�(@���gSQ����:tC��AY[ì� �5�Q�Ȫt��	N�@B��N��8<t- �)<
t%&�} (r3�&�]����93�	C&:p*��/��Z6Ŏ P
��<X6<@	t2<,t1� F:�OL�PrA"�M*� �2II I���W�� 4�.]  ;�t</u�P�G��( �r@�!�X��r+�
.@� VS�>Q�%P� �U3����� c��"Q]:X�"׉6O�!��.� t:r:D���000���[^r ��~PP�E
P�0]�M@W�u_U���]WQ��L������ĉVEX
^_�gSRW��3� ��.� �/6�(�iS&��0.m�@>�	$"���, � Te
<*�
:,4i�29�9HF�]�R
6��LbH�d
 ���T+;L*J�&J�PN� �C Q��R rY_ ,�����PV@a^r[�6V��X*(
D�F3���@m���D�K�0�=u��G�sT��
�a�B� ��@�WU�6!r'�&�t�P ��]�X�VS3�3	
�u	6ļ���I�(��	.=:=' Ӕw:�2		��6 ;�6�b�TU���*R��d�l���rɈ���,P
u)RUQ�P��(�/<�Xw�ظ�*Q���Y�� 
�]Z��c[^ˊ
/2�� ���IX_xG!6����t	
�P6�~6��]X��!��t��.o85�(���hBL+�@ �&;��	IJ0���r
 *u &}�2E �9G�\A  �QUWR��6,�Zs�6_$�]Q#�/a�� rZ�_
�c�U
(Z^]�MY[)A�SR6�L�2N?,� ?w s�Y�l	!2�9t;`2�t� r /��u����-��� �(sUJ���H�	  GIu���WPS�� ��ٰ��u+�K��[ )Z3�-Oa�A�@��Z(U����Z XI)X�B �&�=u�� (��UQ����YU
s٩ȩ;�S�"]q�' �  ��r�ƀ
�u~�>]������W6�>V�&�= �t&:r �:Ew�GG��_�6�`���6�6d���	v���7�0RA2�t<�@u�|
,u6m(]A�$	�a���3��3�Rk�
��!�%� &8%�Qk8e�:�PGK�s �BIu�V���t5M�u,�D� 0�RR<0��74��6�B�>_�uB6IOOEF��W+� h_Ys� Q�H�ʎBtw�#�^��T:	�! :3�#f�nQ
oP@;�DT�|�gH!�tU:C�u�_:'�	2Xg" r`�Y_]^�
���Sr������C[@��y�X6��fC��@A��� ���f"�C��M*1��u3)f -6�	�� ]O� �\�D	:�v*���(]��t
Y�bY�u�I�8Ls*�*`ъ%OC����(�CiB��Wu
��[$[l�7D�X��	`��u���%UÆ(�!˱��>:�[C�5��H��]70u{ PA�B�s�EP�*K etGA��+�D]q L: 93� u&#���u��C$Y�L�u�X�8Qu(&�,����-C{eq.*(U�z,�,�,�@t*PR�82��B�٭�m�
��Z
PX�,���ǈ!	���
�PȲ-RА-| ڃ���"� 4qU�AI�Kn,(��(_(n(�`(4T3�(ҩ�FB:)��@.�▽� �F��f��!-ËD�:=c v�Z�5 @�r��I6:	�Y0 PAAU� ���t�w�  6<|<~
��a/��pj����ti��l�o���i�L�s彚��`@`<|,
�C��"�הY<%ײt;:e.�z���
� ����v��$�������
 �
�t��s�U(������ rZ���((�p4  �P � Z ٘ ,� -  � ./021	 Pl3�4�  Incorrect DOS ve�rsion
suffP(icienmem%�*yNo- (setting syst: &le %1hTidd> (Dis��pla5 M cha�S#+aAQ1ribuMs. 'PATTRIB [+R M | -R]
A
�4A
S
SMI
H
H
[d?�:][pJh�J]Sna�5�/(Q  +�� S�qw�J on-*�C3ar!�
RRd-�only�"$�A"Ar�]΂ vz�.*H5�H*��[/?Process%.i���ll di�o:�.�(�=spi%ed �
B�<)��� #  	  
 $    )  Q  R *i%1
K�	2;�
�	+	, *Co�UgmTeism]�AI� youvu	�T(Y/N)?5PuInv��R��ty� ue���_+�� �(��� Ex�Un`.Err�D%�+��� �$Pt��e!,!�VA���  ���D!N8Df"D <s� �Y� (6 +��� r� ���ׁĎ�s�x�3�� ���L2���6�&2"�Ʊ $��H6���C�@�+��۴J(6�� �����+�C�I�L; ���d3��6�����c�� #� 
Tx.{��yjR���� 5�� ����%��-Y��(�.�y&�, �
Q�#�3۠���s �M6d���N.��.�6"9� t,� � �t�t��3
qJu��D%��� T�����tH���AdJ�����q�r
��P@�t��@Ky��n� 	� �����}ti�^^ fl � �8�#[h�F� ��� � ��_L�^�>q^q��U`)�A� �	���+�(%�>�$�0t���� �;�s
OO������ ����Et������� �	&��{���>�B� ��i�B
�[�Y(P��+��;�r  @���3��E�V3��B 2 
���2�����U���"��,^Ï��B8�,t)�,P
 ��A���3@���u�GDw��Ћѿ;�� A1�]��A�����"GoaJJkGN�)��\X	�=$<\tB��3�A*I���Ӷ�@�Ѩu��91+�N1'�1��1�1��
P���G�� ����+�ģ�����8)bf�6����&���6���ت�O�E !�y��R3���Ji�b�^{'�P����\�J��s)["��.J�4*!�4��64�4�e4͏��  ��&��U�*04���I@B�t��&�>)($ C�E�� E�@$������>W �	 � _����  .���3�I��<;C�t�~ EEq��N�]�Q�V 
3V���;�g@��t���0^���_����W�O��������%���@�!_ )��"r59  s% P�ر���	0��+���Ë��Xr$�HEQ���.2����r\$~�s�6� X� `��2�� �â�c#� >�r<"s r  ���<v���ט
��U�������@�^;��� 	�*�FyH���~o �y�ѸS�&rK
PCFVy(�x,��6�VSއ$$�J�N��V�!JQ��
���=�F� ���E�z�׋ތ؎��*~6�u�A+��GF�A��t�I ������]���@�o��E��xxǨwU3rv$�h3jA�M�^��ґHVW��
�F�͠ �F�<%t
<&t�E�����D�BD�V�'�F� o
�}
 �U�^�]���E
r �v���+���u-Z�s� ��V����PV�b,8�}eS��V�B)�-���,���&&�H���v%v�"����e�`VW��D��!B�� ���=��� H�@�
��]_��Q�׎��t=J^#	^���_��O�W�� 
-CZ\x0da�*� �Ofunct� W-	��5JXMBR;-Time�( Library  4Copyright (c) 1 P988, Microsof�rp "  FILESIZE x (b� D�Ex| � TIM� �U. 
U�?		�Q +A�L-+R2�+S+H�B= " ((&*.2(�6:>=e�i Mj$�Be rN�|�t T �A���-���9	b��K����J 
h �
/�,S�T?  
z����. \Lj�� @��#* 0 Ŧ�sЁ�"b=T��¢e'�P{�		΂<8 n 0�t�
$�N$$�]�0n�p<rN � t �@ ��tS`cHR *.*\ .��.\S����Ar� (	n O[]|<>+=;�)"���V��i]�#$A
!��gV�&= 6 (C) !1-9MB4 *Lcens�M
!at;ial�V�pt��y &/A���Ms��_rv5
R��� Y�L�!�";C_@�>_INFOR��*�-�.CT��" 	�,��("�<<N�G>�BgR60��\ stack�$flow�I3in���g�N�vi)bet�3�k!9!nCQ�ou�UťH��+���.�nm�d.� BY� r�ltleZp�њiE2Exa�[poq��TҶ99'1vlu0#�W�assigc�q����,(�t9 (	2�RB���(D��   	 ��O����P D�4 PˌÌ�H��$� �(l��G��H "�������( +�s*+�����ڶm���� ��¬��N���FF ��<�u�2�<�umm� ͱ�2E!����3ҁ*)����i�����& ���� �t�� ��2[@��)���○>�6 P�� -3��� ��֋����.�/�@	�� �ʨ�q�sN�TP�e�c�is L�$ups 0 �y% >   y � !|"U,�,�,�@�<-�-H=� � �� �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                MZ�   n���    ��R   PKLITE Copr. 1990-92 PKWARE Inc. All Rights Reserved   � * +     ��� J� '                   �>��  ; r�	��!� Not enough memory$-  ��- ���P�� 3�W�D��ː���S��- ڌ͋���������NN��+�+؎Ŏ������ 3���� �+����5����6����;����]����^����_���r���Jt�s�3�3���Jt�����Jt��Ӆ�t��Jt��Ӏ�r��Ju�����.��a��
tu3ۃ�t*��Jt�r#��Jt�����Jt�����Ju����Ӏ�s.��q���V��+��^���Ju����Ӏ�r���Ju����Ӏ�r���Ju����Ӂ�� ��뼬Ȁ� <�u�[���3�����Î����&����Ò���ҋ����S�P�Ŏ�3��؋ȋЋ����� 
      	          	
    :  e r �J� vq
 N�xOb�a���!��?3us7N �4
��,O(�iMl �!Bڦ�y@�y�!9P��07I�m
 �Ԯ!{r���>��$Y �n	ۺ0
����H��tK 7H�t�08!��tK�$��B`u]<�u !]�"#$u]%&'�u()�*M�+n]X,$-�.P./�c�0�15pP� :6��78k� d �<:��nh;�<=��x>n]�?$@�u�A]�F�G�u]lH�IJ�uKNT�OPPTN�0, 25t;4� A.�����.	$
$6MS DOV  ersion 6 (C)Copy right 1981-9 �4 Microsof�@rp LensedQ�at;ial - PR�!pty &Nm/AlM��se2rv54�KSDKHC��. �� �]�A:\*7 /`Z;b�0 hq S����@:�	/V /FiX?�/
�`[]|<>+=;"�I�����~���D�} ? �,, FILE�0CHK1�/\ "i..c. �w�. #K`����
a\�999
`F �ile allocat��ztabbad %PSQR�� ��  $;�~#���
� �! r������+� &�� ZY[X�=V �WU���RP?	� �����%Z]_^K�.ka-hWV'�he��&�,i^_/. �û 3���.؎ԩË�G�`*0�C	�duS�
(�&jC��@��(i���s�������� 0P �W3ɫ3��.�  ��/���>�)m��S��������"����*%(���m��-J
-����@Q
�$$�����
�b��8e�(E��)��. �A Q�P rY_Z  ������PV� c�($!�6Ԃ֪(^�D�\
@3������Dm�K�0=u ���= s�������
 �B� ��fWU�|�� P��t���]$�jVS3�3�u ����%��t�Tļ���U M8=' w�@)Ã���27�����Tͽ��
 � t�T ��� r�u럜+u)�RUQ�P��/<�D�Xu	�ظ�����Y\���( ]Z��b[*^�/W2�� ����IX_wG� ��t=uP�|��lR��  t&�M�	.85u.Q��d-��tP&;�.I%�	I�(��r!�(&}�2�F� G�� �U �WR����6����(N�u�& M �rZ�_P���
Zp@T]Y�@�SA?@�<5,@ 5w s�Y��!�2�6t;��$tR r0����J��-��豩P s��U����H�	� GIu��=  S���ٰ��u+� K��[I3�%L-OA�@��Z�
(UP=�Z �RXX�B .�&�=u�� P��UQ����Y(�s�ȩ;��� "]q�' �  ��e�ƀu ~�>�� � ��@W�>�&�= @�t&:r�:Ew  �GG��_Ï�3ۓ�0�6����	v�(��7�0RA�uP B�t9�u�|
, �u�6�A�"+tuPU�3����e�	 !�%� &8%u
e� t:�uS �s�BIu�V���t3M�>�u+��AD0�<�<0��64��Q�>�GB( 4IOO����W+��
 �_Ys� Q�ʊ�J tu#�*D^��B	�:3�@PdgQ��
m;�D S�|�Z�(t��B��h AT%Te�R\  � rY_]^~
'��Rr������K>P�X���C��@P`��� ���
�"MC��-ۿ$eu� -��� ]  I���D	:�v*�����t
JT|T�u�E (8Ls*T��ъ$����t��ӄA��Uu
�nY#Y؀+B�
�tA J��u�� U�!�z��	ˬ�>9�t�r�KrH$��]60uxP�@A�Z�s�EP��P
�tGA��+�D];�%0��4 r u$"�u��C$8N�u�p�T�u&&���*��+���.�
,(&U��*�*� 	*@t)PR�82���Ҏ� �,��ZX��,���ǈ	����4����-R���s у  u�}� ���6�AF�Y/S* %%X%��g %Zec%0O%u�NB =7J��;,��U�� ���{ �-ËD�)=c v�
�
A�X���I: Uu�0 PAAO��z t�>��q �<|<~�a,����p����t�eT����0��eN��C�v\U\<|,@W
��W��%K�$�8:��_. �-C�	��.hI��|b�����؞�E��r�;��+   B X s �   � � � ��  
 -�E-q  .�/�01C �2�Incorrect��v3��
%1\ �ady ins�)t�ed*�#C$-lo� cha to �f�	(Y@�/N)? UnPo'�K�r%faD dig��QE�[ CB"+}bytR�z(sk space�QQj� As�%2 hidden���vit�u���5�Ұ�C'woul�;be( |aj�vaon-���!mem
�1fEeCaJ4nn$ DSKD netqrU�kA�f)�SUBST{ �pASSIGN�j*&�b}0n-���
�t�uxD�i��g FJ�AT�1+/Ch��kȎ�Rz[	pf��y!tu�*�p;��t..-6(�[�:][[p#(h]na��d]/FV]�w.?  )(QjSppi/��zǻ�v5cL��pE  O�Z�@(s)4%�frag1n��tuF-�66�#�FixB�s��@J.P.݃V.D-�su�wͷ��e�y�OB=;Ty����wiout2vAr:X}s �6cu�+�nt>XJ���:
q? L�[!Uv�����   & 9 a �   �!�"   �# $ 2% X& � k' �( �D�r%1$��%6�A��P�cFguo�b�kscw$�s���d|ʟʷ,PE
Ufnd��, F �Ut� ?�B���oLl �2rwrit/n0 "���cessA��cxXc����&.Vl,e)S	�+>CHD� IRLf�
�4tr�Ryn#�n�! cȹd`�mHa>v�Widq�9X�,�%=H��/I+sub-( ����\o�b��ex�t4��r��;Zru,��= f"A�X /��%sizdju�<M#0�p�:�ܥ�H*p�^Wd��)��i�$�l�m�jpt4JAh�FT�*joBA�frE�ha�f�B��nk	�Bibu��
����
)E*��+ y�x'��$��^ 0 1 D ;5E6 f �7 �8 �: ����< �
�2(5.��{�s�xn��%1: ���=�B,
Tee��th�ptp��gdoQ%;& ��� (r�>d"
��#VLolum�˃Ce%(��%3�!w���sk�� $�<ch*~���=�k���36sP.����.�/�+v�}~�$�#�R�.3	�Àro�A4���%*�O= `�y|��x�C4�q� B *C � D � E ��y� q!H =I O@J4K pL �M$ {N �O 0  P 1Q R 6S Lp�T �!�a��� a<h v	�- #X�[��$suf1i�� �m��� -)B�(MH���fm#�����,oU���		,

�1%4%5��/6���TS��Nb�`ս��>-H�����
[��Ea tEW �&�ault@�8,+D"�,��V�d|*U�9W �ws/DosShea�.Comm��@����MM�� ���Yv�W�㉵i[r꣰*۔*�O�@
oRw�}L�&o��:��A.T�unhQ�,�m�ǘ �+�ՎSba�R2F_�AB67��rac1�D�Vshrēek�;, �MOVy`EV�J�@Eso������-_7E[F�8�,vLm0�N�HELP_�xat�[�fp���"L�tcj�?uT�V����qSCANDI�w� 	��li�P�'ds��c�zfix �muT�wiᲗg�f�˙�ms�/�m�[�)Do�2 you���wt�ac��(�Cv�"��� ��� Ex[�d�)d%9n%�&�� �$tPar�!	��!�U ��� �ڋ�  ]�u�M�u�U	�}8v
�K��]6.� ���b�!.��
�ۋ���  P3��+с� s� �v���K���� @�CP��،�+ظ J)�?R�� ��.; 7Lw�HEZ �	P���X�( ��2<�u�2  �6��
��.��*:�@��Z�ʴT3�6F�G
)�9�E;Nd����?	 �1�G6���G�H��6���H �=�r&�9@b&�:��<�B)>��+&�;O6��:W�R6���J)�	u� ��s	� ��� ��FbU�-%=�P��� ��舽Y�h�  ��G��� P��  ��� ;�s�L 靔$���{�PK۠�����sb�q�� z`��M �u �&�<@=<�t
�� ��L �&��:}�3�PP ��  ����;��?����u� �{o�O�����uX ��s��%�U"�}:u;
 ��6G�5W+�t��ރ�u�PG� �' �_�s���>��(�� �Gc���ӪO�6���)8@�< t&�
:��.���LT�����,AQ
�uYƋv ܲ;>:s$F;x�B@�>�����	�� ��!@���t ��@���r�P�d  �  _F�����6�란���u���JXA#��>BQ7t��%U0���E���2�  ̋�2���HH���� �� ����q���3� �>x���) ��D % ��� ���&�p �`���� ��%�r+������(�����{ BP�}�����ð3ې��@\�f�5�JPr�ږ�� !�uR
(����Z�5ܱq��R�'�_ Ò	8��y�
��\������e�B贠Q� �& @� uOA��r�< � B�| t��.��"O��2�@)�Y���s����@�û.|�
��
\
s���P$��6  �>"�F�_�JR)�JTJ^5��(l��n�7q�v+ej!!&n
!n�: p2�������CU���+s��b$4�bY*+�8�8� ���c)=�#��� �n8��ѝ�O��%� '�Q� ��@ �� ���3۴��r��;�u3�&�  P����ú�"���UcN(+� V��
P����,� J	 C�À��@Z;�tZXUP=�= �S���2����	��[A3�t6v�B�xpQ �0���z��;��y^hz�ƻ�2�Ѫ�.C�A����>9W
� ���&�=�����u��St����ÀRVW�6E�E��ӫ%CWDN6q��C (���^'<_^����3�q�%���q\tQ������&���YXl��ŀW�x���᣾{.��HR�TG�28)�H�9�uPRS�K����Q��m����
���`3�  
�R�a��«Z�5GGW�P�[_[ZX��w������A��FG<�������3�%
�t @�-�/ &�<Y[�/����� �љ C��y�t; >>u
��&��	�
(
F�T�ك>`b�~�5 0u�
�u�� o�RP3�R�x)�`�8%q�χE���j���*SQ�P<R��Ot��� `�Y[�����0�ndֶI�Fes��oVQRN�H���l�
 n$�����;6�p�MW|�r5w ����u^���.�v���"�`eK%�.JTKK_�	(e�C ��ZY^B���� ��v��+P�|2�*�15 �3�`-P���=�t���5�B ��TeX_^e/e�Y,�2
#	;�)� V.�@;���߳XX)b(
���Mx|R����6SS_6dE[W6��O(������z�(�QP ��RQW�-�s�PXP��2䣀�� ��B�XY_Z�����Y:
��-x���.�"�F���.��jx ���J�����m��#N8	[���:	|<Y	>+H(X	=;K ����S&�&:s  � [��6�SWU�  ��� u>��rr7@9��t2��!��� AtN��<=�PC�^sɬP C��NP�� ���j�6W�</t�Y1"t>�	��G�P�9�s�@��CC�-� �S9f�^U
%@�ăk�CS�(&��s?3����++3U�+
	@�5T5
5 ]�_[�?���������� 2��� u���u��uBg�P� ^��� XƀbX���UQiO j�o	�)s� �@����.�SY]�&��`~ �E��E� �1���rB�& �
�P��+��XlD��r#�|�
�s	s&
��?<&��,�g�-� c��
���0�Z$ʃTe[~&�EX�G<C�ULM�Y<u H�O<t�<t�<	��=<u��@,J7.�].+� 
u
P&�G~e��&	�t�&�-Xt5D_��A�AB���WĄ����_����<�� � @����>V�)�X�S}� t	� �>*�d� x'saX�PVbt<:`u�|*� @'�sFF��^"�R��A�L�r*� �� ��Z^�<�s  <ar9<zw5$��1SW@�>3	8t�QR�De��I�e4VO  ZYX�]�ECC,�&�_
�[B0r<9w,0���X��u�����T�@�%URV�T0� �:�{�!t��W2�n���t�
HAFuZ�Z&:FI�	�PFE#�lCFHE
i9�7@t&�D>G Z(ȁ"E ��%	M�7P:�t�����^Z]�WV�>��W�W&  ��^���9]�-�%X "��*
��LsGF��$���.G�>�^_X �	P(��M�gSQ�8	�	?�Q�(�AY[{RI5�@9r*�|�- ��   ��,`\��K���T$ZT����R�Q+��t�	N
$%��N��x<Dt-�)<
tQ %r3�@�&�]��9HA�3�	C&:�����/��6�� � ��<X6<	t2<,t1u��� F:��P2	�AM%����2II Ip�2	A 4�. �;�t
</u�̭��
@� �VS�>��%`DPQRWU�  ޸ c�!���]_ZY�Xȉ6��(�����:�@r:Dw�����[^ ��o�[1��
 }莐_�t$�N��
q8�r�
���	��(�����
D���R-/*����LP� ��ي\  �	q���� ��"��ˊ�b �{'���(��W� AA�x�� ��0��U&�ک��K ^�� �>m
�� &(�	�&:�tG���&�E {��3�3ҍ6"&P�@�V��=��DBA=
�; ��N"��Q<*wN���DBM   u�F�6� k�ܣb��-�����-Pma�u!E �&h�ύ���>�P�u �F���2t��{��Xe*V�K(z(e�
8�2m }�L7 tC��t�Dt �6u��&��������`�_Y�縀���w�(֜"���"���2$�� T���*��� u�@=���c	�s:g>��^�ѭ��P!`$�E	e��+��s(��(O��GF4�������sE���E� �%J��e�C	S ��)��ËO�QDɊO���Ht���T3��DEG	=�%=�( ==i�t=e=�0>=@7� =�3��Gt���SRP��5� �$G��[Z�@�o��т	[G
i
�(�k
�g�6,�hS�[D�	S3��2�ן��'�E5�,�, �0�� t�貧���t�唲�Å��2:*��2�AM�� �X!�6�ȝ'�`PB�#�5q��E����>���%(�$�V��ʟ$� D[�
 ���/���������  *����T�5��u&(W� (��t0�C I�
��[4���T��F$ 0ܵD�E�S�Q�+6�t�5� ��WV3�3���@��������r��@��s�r�Ƌ��03�3�^_Î^�& ��&I;uG� �c @��u&�=oxu�&�}G�Ã>�R �3ɶ�@�� �ոSJ��դQ�����r	�:��NuxEQ �VR���@���% �^�龋Ha��茰#��e��0Zr\��^�2�Ck ��j�����(�p)�[I�p�o P�$��:dt>�@�!�'��'G��:����t�� �(MO�L&H�W룴��֛��Caj�	�+S6������n������
�3�-%P�(M�X� 
D��V����9~�0E^! ;�����t!�s��@a�8��pu�2��� ��YË6-T��>��]t�����5q�RH�T"�
 ���6�t�:\ҍ���7�_RV�� ��)���Ξv��W8�����uP��X�@"X.���NXX��`m
��o�.�B���.�BR4�ȴM�� �1�P�'�˴,������
΋�R�* ��������
�P����Z���EP&���tA�� ��&% J&�6���&��ȣX&�6��A��䀰����X�8к�ֵ5�U������� �N��3�S`�U�]U�qK��,�r�P-3��� <����
R��(�+�F
Z�<��ZXo�z V>��][X��f�v=va���v���	(wwu>�:�d��d�d;d�&By �,���/�t���U/6t~������� 0��v����A���]�
W
s  9 U���,;&w����k]5- �����w�| 1��W�,�Z���i�~|���*�!��ss@l7�}��������5��]�p ��X�j�t �P��sX�H��X���D�uVP ���9��^�L l��D";Ft�������$M	�&��b"�"��"3�!$&
c�c$ӴV�*t��?�����v}�}^cc}&V~t�i}D}��}
}	}Hve>�� ��+:tȁ�su(nu�*8p����1�,TY����w �tu��N;�7	F�m�5  �ڠ����|PJz>>&<�b���5*�Qȃ Y�"D$�2 �M��Bw�q5��ƘDg1&fs��T\33�H%Z.���.�d���AJ@ �6S@P��@v���L3,�X_� �=��r X�e�[��AND�u4�b���`��8 ��Dsu��������!?&��� u����b�"M��T�6U���Gpz �PW���  �^V�t"�<�^[]`	�T&*�
�1�I�v�B�Bp.j��މ��ދw2�k�uSS��[�'d���t��?�6/[AO;�vD�!QWx�6hK���:) 2w2Y�#��t�8 ��~�6#�3��K���9��GE *�$�>�78 2��&��P���+G b$W&r
�u�rRZQ�w��&�F �PfJY���Y�������ZR� Z�B�3�2�+".w.�!N��QJ1�$j�&���y�VSQ?���Y[^��USVV`\h ^ �c���l�  `Ë^;:r���? �������uR��s�(���6ՊȤyj�j�P�����ަ��w�c��&A�st�X����^��@���Z�÷���`;����t�%
�c��V��w��y�^V�J ]@��:������/>e(	F�i�N��^��8EG	`�t���� ������C�F�r�@>y:\u�{E)ܠ:x�t_VS"��0��aS�C����x��9��AAT>T�Z�|"(�$l �
Pg�;�8�P��&`n	�Xs'D���u=3SV����A�OT�^[P&'��/�[����p^��d�v��� o	�r��"IVW�SMȂ��[_1�tW���D_u'A�t[����D�J ��
$(�GD&
��:�������<qg�m�Z��LVP�_A�X#��d�߸v14�1yA	@�Bt@�Bu;�s�>�3��
3)S@+�Ӄ��
/'>r�� �X�P����� (���[�P�Xy�X4
�����<�^[X�V�����4m �&�ּ,�27 ��    % 0 ; F Q \ g � � � � � � � � � � � 7���Jf�(F)�)�)*.*�192G2�2 3 44T4�4�4�4 �   '                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               MZg    22� 0fY       �&  �    k!                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              U�� ��F�  �^�������P�[[�F��~�|� P�[��]�U���R����P�v�[[����P��Q�[[�t����P��P��[[�u� �>� u�v�hP�%[[�v�[� �����t��v�)[<u�v�0��v�P��[[ǆ��  ���؉^����t�G �F��~�u&����yt����nu��P�[�~�u:����yu3�z��~�t*�~�t$�~�yt�~�nu��v���[� P��[�F�����돋�]�U���TWV�o�^�7�P�$[
�tl��P�DP�[[�t��P�^�@P��[[�u�� �3��P�^�@P��[[�u�m�+���^�@P��P�[[� P�[�N�F�~ u��~ u�xP��[� P��[�F�  �p����P��Q�y[[�t����P��P�g[[�u"�^���v�0����P�[[��P����P����^���v�0����P��[[�E P� P����P� ���F��F9F�}2����P�^���v�0���|[[�t�k�����P��4��P����+�P�7[^_��]�U���V�^�Gu!�Gt�G$��P�v�e[[�ub�v��Y��P�� P���[[�tE��PV�[[�t7�v�[F�F���P�v��[[��P� P�v�X���^�� �v� [^��]�U�츠P� P�v�2��]� U���>V�>��t��� �F�n�F�5�F�P�[�F�P�N�Q�N�Q�/���F�F�FЉF�+��F�^�&�@��B�F��
|�+��O�B��=D uE�B���؉^����t-  ��B��=N u'�B���؉^����t-  ��B��=P u	��
u+��&F��
}�B���؉^����t�-  뛊B���j�*����^��]�U����F� z�F�  �F�P�N�Q�/ Q����~��u� �+���]Ã>��t�����Hu+��������u� ��U���
�, P�D[�F��u+��EP�v�v����t	�v��S[�Ḡ	P�v�?[[��P��	P�[[�t� ��	P�v�~[[��	P�[��Ƈ�	 ��	P�[�؊��	P�s[
�t��	P�[= v��	P�[��Ƈ�	 ��	P� [<u,��	P�q[= v�^��.t��Hu��P�s
[� P�	[�P�D[�F��u
�v���[�7�P�v�3[[�v��#[F�P�v�[[�v��[F��F�F� P�v�
[[�F
P�v��v��V���v��0[�t��v��e[�v��0
[�v��)
[� ��]� U����F� C�F�F��F�PP�o[[�~� t�����F���]� U��V�^�? u�vS�#
[[�E�? tS�t
[�^���@�P�5 [
�u�(P�v�	[[��F�^�P� [
�u��v�v�	�^��]� U��~\t�~/u�]�*�]�U��~/t�~-u�]�*�]�U����F�  �����F��^�P��[
�t�^�GP��[
�u,�v��v�� [[�u�v��v�� [[�t�N��v��	[F��v��v�([[�u�v��v�[[�t�N��v��	[F��F�P�v�k[[�u�v��v�\[[�t�N��*P�v��#	[[�t=�,P�v��	[[�t-�v��3	[F��F�P�v�� [[�u�v��v�� [[�t�N�����P�v�[[�F���]�U��V�^�? t�:u��v��G�D�D � ��^� +�^��]�U����2P�v�k[[�؀? u�F���@�F����]�U����*�P�v�(
[[�F��u�v�y[F��*�P�F��F@P�
[[�F��u�F��]�U��V�*P�v��[��V�[[�t�,PV�[[�u�6�V��[��V�v�[[�^�?�@^��]�U��WV�*P�v�5�[��W��[[�t�,PW�[[�uW��[����W�5�[��W�v�f[[��+�^� �^�?�@^_��]�U���v�v��[[�t�v�[F�v�v�1�[[� �+���]�U��WV�^�? t
�:u�F�v��[���v�v��[[��+^�~� �=�@^_��]� �9
�u����!t�8���9���À>9 t
�9 �8���!2�� U����F��F�F��N�QQ�[[�F�N�F�F��F�F��F�PP�[[�~� u�F P�[�F���]�U����F��F�F��N�QQ�b[[�F�O�F�PP�T[[�~� u�F P�F[�F���]�� U����F�C�F�F��F�F��F�PP�[[�F���]�U���WV�F�F��v�< t�|:u�������t� FF�P���[
�t�DP���[
�ux�F� �^�? t*�:u$���؉^����t�F�, ��^�,@�F��F�F�P�v�[[�t� �l�F�^�?.u#� t�GP�o�[
�t�^� u+��@�v�^�P�P�[
�t�v�v��0�v�l[��^�G��F�P�*�[
�u�:P�v�[[�v�v�[[�~�~�^�? u�� �<P��V�� [[����F�� G�?PV��[[�u�F�N9Fs�<��^�P���[
�t��[�APV�[[�u:�F�N9Fs���^�P��[
�t�F�N9Fs����^�P�y�[
�t��V�v�?[[�v�[F�F�P�X�[
�t�F�\�F��^�F�
�t�5��v��i[= u�^��G\�G �v��� [��^_��]�U���v�v�$[[F��]�U���v�v�i[[F��]�U����~ u�F��F�PP��[[�F����F�F`�^�F��^�F�:�/P���[
�t�^�F�\�	�^�F�/�F�G�F�F��F�F��N�QQ�u[[�~� u	�v�k[��� �F���]� U���v�Q[��]ô0�!<s3�P˿�6 +��� r� ��ׁĮ
�s�:3�P���L�!�Ʊ��H6�J�L6����6�g���P6�g
��P6�g6�g6�&F��6 ��+��۴J�!6�������
+�3���������3��H �6��6��6��x�P��.���ظ 6�H�P��6�>���uXP6���� P�H � 5�!�r�t� %���!�>� t6������&�6, ����3�6��s�Y6���ڻ 6����&�, �>��3�&�= t4� �d�t��3��u!��������,Ar����,Ar
ª��� ����� D�!r
�t���@Ky羴���� ����� �U��3��U�� �U��VW� �U��VW�Q
�u����� �����v �>���u�������a �����g �}�tX
�Pu�~ u�F� � X
�u�F�L�!_^]Ë��� ���r� %�!�>� t�����%�!�;�s
OO��������;�s���Et�����Y��+�r
;�r����Q3��)� U���WV��V�������FP�v��P�p���F���PW����F�^_��]��J �% U��׋ތ؎��~3�����u��~������+����F�� t�I�������]� U��׋ދv���؎�3������ы~�Ǩt�I�������]�U��׋ތ؎��v�~3�������+��t������]� U��׌؎��~3�������I���]� �����
�u������>���u	S�����[��!� �U��VW��
�F�͋F�F�<%t
<&t�F����F���F�D�F�D�V�F��F�~��]�M�U�u�}
U�^�]�W�~��]�M�U�u�E
r3���� ��u��
_^��]�U��VW�~��]�M�U�u�}
�!W�~��]�M�U�u�E
r3���� ��u_^��]� U��VW�~��]�M�U�u�u
�~��]_�!W�׎ߋ~��E�~��]�M�U�u�E
r3���_� ��u_^��]� U��^�_��O�W��]� U��V��>���u������!�� ]�U��W�~��3�����A�يF���O8t3���_��]�U��^���,A<sa�C�
�u�]�U��� VW�v�Ў�� 3��~��
�t���Ȱ������C���v���C�%� t���Ȱ������"C�t�_^��]�U��� VW�v�Ў�� 3��~��
�t���Ȱ������C���v���C�%� t���Ȱ������"C�u�_^��]�U��9�U��;�V�!��U��:�V�!s�= u쒓�C< t
<?t<*u�����U��V�A�!� U��� P�u�>� t���� P�c��]ø �:�V3��B 2���2�����Ut���� P�<� ^Ï��0�!��� <t)��&�, ��3��� �3��u�GG�>������ыѿ �� ���< t�<	t�<to
�tkGN�< t�<	t�<t\
�tX<"t$<\tB��3�A�<\t�<"t��Ӌ���Ѩu��N�<t+
�t'<"t�<\tB��3�A�<\t�<"t��ۋ���Ѩu���>��G���B���+�ģ����6�?CC�6���
�u�6���� �3���< t�<	t�<t|
�tx6�?CCN�< t�<	t�<tb
�t^<"t'<\t���3�A�<\t�<"t�\��Ѱ\���s�"���N�<t.
�t*<"t�<\t���3�A�<\t�<"t�\��ٰ\���s��"���3���  �&�U����&�, ��3�3�3�����t&�>   t�F�u���@$�F����	 ��P�������ϋ�3�_I�&�6;duQVW�d� �_^Yt&�?CC��
�u���&�]� U��VW�V���;�t@�t�3��������_^��]� U��W�v����t ���3�������I� �>���u���@�!_��]� r3���]�s�P� X2��]�s� ������]�2�� â�
�u"�>�r<"s< r��<v���ט��Ê��� U��VW�v����t����t	����uH�������v�Du8�u3��t�D��D �E �L�� �S� P�	�[[�t���3�_^]�U��VW�v�������v�t#3ۊ\���@tV�LX�~ t3���E��D_^]� ����'P�U��q�M�VW3��F��F��v��v�F�
�t�~� }�F���, <Xw�$�� ���F������F������.��:�V�� �#�3��F��F��F�F�H�F�랊F�<-u�N��<+u�N��< u�N��|�<#u�N���q��N��j��N���*u�V�y�؀N����02�F��
 ����F��>��F�  �6��N���*u�"�y������02�F��
 ����F����F�<lu�N��"<Fu�N� �<Nu�N��<Lu�N���N�����F�<du�<iu�<uu�<Xu�<xu�<ou�<ct<st'<ntQ<pt`<Et<Gt� � ������O� ����u���u�w�}��W�N��2��uOY+�����Y�F���F�t3���>��F�0u�,�9�/�F�u0�F�� R3ҍ���� �� ����X3Ҿ �Ɔ��:�	 ��F�� 3ҍ���� �p� �����G�F�N�@�F� ����~� t�F� �
=g u�F� �����v��v�VW�v�F�t
���F
����F��
�F��t�~� uW������gu�F�� uW����&�=-uG�N����W� �OY+���� �N�@�F�
�5�F���F�'�F��t�F� �F�0�QV��V��F���F��t�N��F��F�t�� ��� �F�@t��3��F�@t�}�N��؃� �ڃ~� }�F� ��f�����u�F�  �~��N�2�v��5�F�t�&�=0tO&�0A� �F�@t1�F�t�F�-�F� � �F�t�F�+�F� ��F�t	�F� �F� �F�+�+F�}3�WQ�F�u�Ȳ � P�~�N�� X�F�t�F�u�Ȳ0� Y_P�k X�F�t�Ȳ �{ �	��v��vËv��Э��v��F� t������������u���ØW�^�Ox
�?��3�_�QRSP�� ��ZY=��u������N�W3�&��������_t�F�����N�W3���������_t�F�����W��
�u�u��3������0<9vF����N��Y+�G��_^��]� U��V�^�L9\sKK�9\v�\^��]�U��VW�N���w�L��s�Ur��s3��� _^]� SQ� ��QP�{�[��Y���t[Ë��S� U��VW�v�D��th�@ud�D  �t�tW�L�$�$�D�������v3ۊ\�uL�u�uC���t���t���u$���@t� Q�~WS�k��� �>����L �\SV�[[�Dt֋�T+�B��UJ�T� QQ�tS�1��Y�|�V�;�u�3��F�3���� t� QPPS���3�����_^]�U���WV+�9~u	+�P�e �U��v�D��$<u:��u�ށ����vt(�+D�F��~P�t�L*�Q���9F�t�L ����D��D  ��^_��]ø P� �U���WV��+��~���F�����96r�D�t�V�\���@t�G�䐃~u����F�^_��]� �A���S��w�_
3��#��[�uBS�w�_;�t6K3����T�;�s��r#��t���H;�s#�r�Э�t�� ���D����[�G�G��[�L�t	�+�H�+����ƌ���QW�Gtc�� ����t+�IAA�w�tL�s	3�����0�?&��=  t� �;�r��u��"��r���H���s3���#�R�. Zs���t� ������+W�G��w
J�B�����w
_YË��GtJ�wN;�r9W�s6BSQ�ގƱ��u� �Gt
Ƌ�+ÎËشJ�!Y[r���GtJ�W�����W�w;w
u�w�=��t��$����OO��_� U��V�v� P�:�Y�ށ����v�t�L�G ��L�G �G��D�D  ^]� U����^;�r� 	�*�F �tH�~
 t3ɋѸB�!rK�F
 uFVy(� ��6�V��F��ѸB�!FVy�N��V�� B�!�؋V�N�F
�B�!r�������U����^;�r� 	�����>���u����� t�B3ɋ��!r�����tn�V3��F��F��WV����f��N�8�
�uJ�� =� vF���ܺ =(s�� +�ԋ��N�<
t;�t����" �j�;�u� ��
�F���� ��^_�^�����PSQ��+��Q�^�@�!YrF�;�wY[X��ß���~� u�s�	����@t�^�?u���� ��F�+F��f�^_���N�u�����V�@�!s�	���u����@t
�ڀ?u����� �� Y��;�s+�����3���                              MS Run-Time Library - Copyright (c) 1990, Microsoft Corp Deletes a directory and all the subdirectories and files in it.  To Delete one or more files and directories: DELTREE [/Y] [drive:]path [[drive:]path[...]]    /Y              Suppresses prompting to confirm you want to delete                   the subdirectory.   [drive:]path    Specifies the name of the directory you want to delete.  Note: Use DELTREE cautiously. Every file and subdirectory within the specified directory will be deleted. %s
  B � � � � � $H���Delete file "%s"? [yn]  Delete directory "%s" and all its subdirectories? [yn]  Deleting %s...
 Required parameter missing
 Invalid switch - %s
 .. . 
 y Y ? *.* .. . *.* . .. *.*  ����*.* 
Deltree has found an error in your directory structure. Run ScanDisk to repair.
 \ . ..  : \/:     \ \/ . .. �  �                         _C_FILE_INFO=                             ���                     �         ���          (((((                  H����������������������                                                                                                                                  ��     	���  �                   �                                                                                                                                                                                                                                                                                            n             EEE50 P      0PX 000WP         ``````  ppxxxx        (null)      ������          ���                  �<<NMSG>>  R6000
- stack overflow
  R6003
- integer divide by 0
 	 R6009
- not enough space for environment
 � 
 � run-time error   R6002
- floating-point support not loaded
  R6001
- null pointer assignment
 ���                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                MZ^ � � @   ��1 ��  �@                                    � A ��   �   �   �   * e������������������������������������������
������"�:��������'�F�K��������� �4�H�_����������6�O����������� �R"�u)��)��)�b*�g*��+��+��+��+�D��H��S��S��U�)V�9[�d[��  �  ��I��c��k��Ղ�奥��D��I��Z��k��|��������������Ѧ�⦥���.��3��ݧ�;��Z��ݩ������%��e���������  �             e�e�e�e�ee�enee{e�e�e�e{e�eD��e�  ���Ӱ�尥F0e�0e�  �� �� ^  B  Ա�ֱ�ܱ�ޱ�䱥汥챥��������������������������$��,��.��4��6��R��h��ڲ��7eCGe�He�  
� �� �� �Xe1[e�� �� 
  �����$��L��Y���
  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
  �� �� �� �� 	� X� k� �� �� �� �� �� B� �� �� �� K� ݷ�ⷥ�����&��.�����                    ��   �L ~ EMMXXXX0� MICROSOFT EXPANDED MEMORY MANAGER 386���   �L ~ $MMXXXX0.�.�
W� ���&�>��3Cu.�� u� ����=�u���_�.�.�
             1
EMM386/Windows interface failure.  EMM386 will remain off.
$                 %  �  fS�  �ۀ�s3ۊ���.��� f[˴���2��� u��>�u���< u�� �
 E�c<u(�>��� �>� �� .�>	�� ���
 $�Z<u{�����>�u.�>	t�>� � �&���
 E�>� t#�� u>�r���2�&�����
 $�� t�&��P���愰 �� �X�>�u ����S< u� 	� <uK� 	t?��
rf��   u��
r(� 	���� u�>�u
��r
���  �T���l<uc� 	t���
rf��   t��
rـ& 	��&���>�u�>� u�&�����愰 �� �� �� t��� 愰慝� �[˴�� ���     ��.��
�ϸ�V�g�                             )            fPSfQ.��  �� �Erz �f%�  .f�"ذ��pf.�f.� �f  �"��:� �(  �3� �f3�"ы܌Ѹ ��f���� f���� �.� �� �Ћ� �p�� �؎������fY[fX���z�fPS� ��&�&- ����z�ظP �؎��Ў��谀�p �f%���"���  .8	 �"؎Ӹ  �؎����� �p�&����[fX�PSQ�X%�P�����؋�j h  j h  j h  j h  j Sj Qjh 0j h  j h)fσ�f��   t��  u� Y[Xô�.f��   t��b��.f��   t��P.f��   u�P u=���d.f��   u�; u(���`.f��   u�& u���d.f��   u� ��R.��
Z�t����Q+��d$��Y�           p �.�� �!��    h� �& � .�.�P��.��@.f���   �愰 �� �X�            .�� t.�.�
.�.�                       �����t+���tJ���tY.��u�.�.�.�&��.�� t��z���.�� t�.����U��P�X�F% 	FX]ϝU���  �ء��f�]�.f��   t�.f��   u�.���fPV&�?w)�6P&f�.f�&f�G.f�D&�G.�D�ތΎ�&�g�^fX�� �.�� t	.�&�����f3���&f��.�.�s�<St<Ru����                ��6H � �e�&��� ��f�^f��&�� f��&�� &�>� �^�� ���F��&��F��&��F��&�f��g�$��&��F e���Fe���F$e���F(e��e��� e����faf]e��e�&���e��e��e�&�e�.�����.�.�
        � �`���� ���r�5H ������aÝ���PSWV���.�� S�h  ��
[�u.�&�߸ ���&�>��3Cu.f��   u���u���^_[X�.��@ �1 QSP3�3���� A3ہ� w�.��
�u�Q�{���[.��
X[Y�.��@ �3 PQS3��n�A�� � �.��
�u�.�>�
 �
 .��
�6���[YX�� �؀���G������ ��             [   `�p�H� � J.�@a��h�            �	                                                                                    @                                    �                 ��       ���                                                                                             MICROSOFT           EMM386 4.49           �	�	S�����s�.���	[�.f�&�����.�� �2 �.��� �!.��`f`.�>�
�Ǎ>�
 .��
fa� .�
 $����.�� �� .�&��� .��.�&�h� �& �-�������rYjPh� �e��e�&�jXe�&��sXH e��e�&�r�5H ��r$.��.�
 E��!�.�
 $.�&���� �	�!.�&����.��.�&������P���愰 �� �X�                        �� g� T� �� �� .� S� �� �� �� �� i� �� ���.�.�
��.�.�
�����(�<������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������
EMM386 Privileged operation error #xx -
Deactivate EMM386 and Continue (C) or reBoot (B) (C or B) ? $
EMM386: Unrecoverable privileged operation error #xx - press ENTER to reboot$
EMM386 has detected error #xx in an application
at memory address xxxx:xxxx. To minimize the chance
of data loss, EMM386 has halted your computer.
For more information, see the README.TXT file.

To restart your computer, press ENTER.$
EMM386 DMA buffer is too small.  Add D=nn  parameter and reboot.$
EMM386: DMA mode not supported.  Press ENTER to reboot.$xxx
EMM386: Unable to start Enhanced Mode Windows due to base memory back fill.
$
EMM386: Unable to start Enhanced Mode Windows due to invalid path 
        specification for EMM386.
$                                     jPh� �h0�=  u�>  �u
e�>	� � e��e��� ��f�^d��f��&�� f��&�� &�>� �^e�>� u �� ���F��&��F��&��F��&�f��F d���Fd���F$d���F(d���Fd���Fd��d��� ��f3ۻ� f��&�� f��&�� &�>� � �� �Ћ��� f`h  �Ȏ�&��&��&��UP䡢�!�� ��!���p�u�X=  u�  �g �% �0�.�[= u�� ���)G���"�� �� �� �1= u���B ������ �%�= u���9 �%�	�h �N �� ����؎���� ���� �� ������ t�:t(:u�@ ���r   ���p� � �q�� ���d��� ��2����桠�!� �p]fa�愰 �� .��.��.�&�.�.�.��.�&��PQR3ҹ
 ��0���0�UZYX�PQR�
 3����tR���Z��0�GZYX�0123456789ABCDEFPSQR��б�������d�G��}�ZY[X�           �d�t� ���d�`<s<��� �P� ���dX��Q3��d���Y�%Y[<wr����f�f`f��f���� �� ��f��g.�E�  faf�g�E�Ü��OQH f��f��ef��e+�e+�f��E�gf�Mg�E á�+�+���+����� f�6�f�>�;�t&g�,�����
shN;�u�f�6�;6�vz� f�>�)�)�;��5 ���f��gf�4�����gf�<������gf&�g�� f3�gf�~��gf�g�f��&g������ ��&gf������% �gf�Eg�E �g�E�����- ��+�� �������OH �V�����|� ��OH ���A���� ��f�6�f�>�;�tN�� ���g&gf������%��f;�tN;�u��-N&g�$�    �����g�E f��s����OH ����g�E������pf��gf�D$ 0 �� �� �f�	f3�"� �f%�  f	"�f$	f,	 4	 6	� �pfϰ��pf�n h � �� ��f$	f,	 4	 6	 �% �f�	f�	"и �؀&- ��� ��fS �f%�  gf��� �f�"�gf�Fgf�@gf�^���g�d�f[gf�Ffggf�Ffgg Vg ^j g�vgf�v� �pf�����p�� ��X���jfU���lf�&nfrfx ~ � �f�` �% �f�df3�"� �f%�  f	"�f$	f,	 4	 6	�<	(�P �ظ� ��3���� ���f�&�f��(f��f3�f�F$f�F f�Ff�Fe��f�F��f�Ff�F 0 � �pe�&�����pXe��ef�`"и �؀&- ��� �� �f%�  efd"�ferfexef�tef�����g�d�e ~e �e�.he�lef�&n�� �� ����f]� �p�&�� �f3ۃ��&g��     �� &g��    �� &g��    �� &g��    �� &gf��    ;6�tiruf��+�v����f��f����gf&�g��� f3�f�>����gf�g�f��f�>���gf�g�f   gf�g�f   gf�g�f   gf�g�����f�����   ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                �� SQRVW�  ��3�� j S���
[=$ rFP��� f��@gf�E   - r���
�X������;�s;�t��S�	��
[�tROu�Z�t�
��
���_^ZY[��b �  ��S���
[;�s=$ s�.��P�д	��
�tR���
�t��f����ZX�Z�
��
X3��� �  �ش��
�
��
�U���F	t�]�                                                                                                                                                                                                                  ���uHh  <tE<u:f�&������b	 �>�t$�
 E� X�>	�t�>	 u�
 $�� Q�.�.��� u'�>�t���
r3f�� �  u!�� u5�
 $�́� v��
 E� Q�R�(�R�xP�Ȏش	�!XZ� ��
 E� X��.��P�  �ظ ���� �!X�       �e�� t	e���g�e�>�u���e��e�&�h� �& ���i� �� e��e���  �  �� jPh� �h� e��e�&�jXe�&�e�6�e�6��&K���t�P7H ��h<H e��e�&��� u�>K@t�5H ��
� e�� e�����
� ��e��e�&��e��e�
 $e�&������������������     .��.���PSQRVW�.���G<s��ྎ�.�.�����G_^ZY[X˰�����3���.�>� �
 .������B�g��PV�&�.:� �����.��3�^Xð���G  �� u&�% &�E� &�E  3�ð���G  �P��  ��ue�� &��Xð���G  ��P�h  ��u�e��&�e��&�E��P�h  ��u�e��&��� ��&�Ee��&�E�fS�h  ��u!ef��f��   &f�e�b	��&�]�f[ð���G  �� ����                        ��?t��t��t��
t��t	�fZ.�.*fRf���   ��r����
s�.f�s���� .g:�  v��
.g:�   v�fZfSfQfRfV�h  �d������.�*�rd�� u�.��d�&����f^fZfYf[�     U���h  ����u'h  �{ td�����KP�X�F% 	FX]�df��   tj@�{ u.�>� �t.�>� �t.f�>� t	��].�.���]���ރ�f���ހK�r f�w&f��f���ۃ�V�t����U V��f�f���3 f��f��f��f��f�f��  
 � f���G����I�" f����^;��	 f�����^f�Df3�f��˃���VSRQP�6B�  � 3ɸ l�!� �ش>�!�XYZ[^�    j�������aaaaaaaa�������fQh  &�� t��sf��gg.�$M  fY�.�.&f�>�   t�fY�.�� �#&f�>�   t��&�>� t��&��@�!fY��PR��  �����d��
�tdf����ZX����P��  ��d��
�tdf�&����X����P��  ��df�&��� C�/<�u!SR�C�/d��
d��
df���Z[�X���X�        .�./�.�3f%����h  �d�� td� 	tf  � ��P� X� ����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               ��   �  ��   �  ��   �  ��   �  ��   �  ��   �  �   �  ��  �  ��   �  ��   �  ��   �  �  �  �? ��  ��  
�  ��  �  ��   �� ��      ��      ��      ��      ��      ��      ��   �  ��   �  ��   �  ��   �  ��   �  ��   �  ��   �  ��   �  ��   �  ��   �  ��   �  ��   �  ��   �  ��   �  ��   �  ��   �  ��   �  ��   �  ��      ��      ��      ��      ��      ��              � H  �  � H  �  � H  �  H  �  4H  �  IH  �  fH  �  �H  �  �H  �  �H  �  H  �  ,H  �  BH  �  XH  �  zH  �  �H  �  �H  �   H  �          �H  �          �0H  �                                                                                                                          �H  �  �H  �                          �H  �                                  �H  �                          �H  �                                                                                                                                                                                          %H  �                                                                                                                                  �H  �                                                                                    H  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          ��   �  ��   �  ��   �  ��   �                                                         ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             � H  �  �� �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 ����                                                                                  � � � *!�!1"8#D#�#�#!$k$�$�                                                                                                                                                           ��                                                        @ @       �               ���          �        



 ��� ��؇��� ���  ��� ����	�
�����؇���  ���  ���
�
��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        �  ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������             ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������              @ �                                                                                                                                                                                                                                                                                                                                                                                                                                                              fU�P �ݽ� �� ��e�.���rB��VtH��e�.��  f����&f;.�u.f���F t��v�v���t&�P7H ��f]f�e�.�f����f��e�&��jg���h<H ��f]f�           fUf���F tj ���  � �(fUf���Dr�F tj��� � �(f]f�fUf���F tj��~Hu�~�2r
�~	3w��2�nrf]f�jfSfV�� �  ��f��f���j j fUf�� � �(j j fUf�� � �(fUf���F tj�5� � �(j j fUf���F �� � �(fUf���F tj��� � �(�ۇۇۇۇۇۇېfUf��jfSfV�� �  ��f��f����
� � �(fUf��j	fSfV�� �  ��f��f��gf��H	  gƃL  �
�	 � �(fUf��j
�� �
 � �(fUf��j�� � � �(fUf��j�� � � �(fUf��j� ���F �!� � �(fUf��jfSfV�� �  ��f��f�� �f��
f^f[���$rf]��fϻ � �(fUf��jfSfV�� �  ��f��f����	� � �(j j fUf�� � �(fUf�� � �(fSfV�� �  P��f��f��gf��H	  gf���  ��,;�tX�x	f�^���.g�]]  �^�Xf^f[��!7Mf��P�a� � �a� � � $��a�a��u�X����  �F���+1.�������X
�����������������������
�������{
����	����
��������
��������������������������������������
�
�������
�
-l��������������������������������������������������������������������������������������������9�G���������������������q�������P`��

�

 �����������fSfV� �ۋ^���� �^���>� �^���� �^���>� �P ��&�   �� �ۋv�� ��.�������h� V˃�V�n�� �ۋv�^�f���\�^�\[��� �ފ_�2����8 ��f�7�vf���vf^f[f]��f�&�  F�v�x&�  ��F�vS3��N&s�[��F�vS3��>&�s�[�SR�T2����v3��%&s�Z[�SR�T2����v3��&�s�Z[�F�vSR� ��%s�Z[�v�F�vS� ��%s�[�d�SR�T2����v� ��%s�Z[�I�SR�T2����v� �%s�Z[�.�F�v�F th� f�� @  f^f[f]��fU���������&�  t	F�v�����&�  u�]RP&� �� ��F�����8��0t��u� �!�  �F�v�߀���� ���&�@���&�A��t�����@t���u�&�A���v�
�&�AF�v�ߋF ��� ��|-t��t!|9��@|t�F(�-�F$�(�� ���@�� ���9�F���ǀ�Ft����t݀�t�S� �Ë���&�� ��&�>� �� ��[U��v�^�n>� ���FU���t>��u�F�4��u�F�*��u�F� ��u�F���u�F$����&�>�� �� �]XZ��XZ�^f^f[f`�^�  �(�.�&�  �?fP�� �Ê&�l	F������&�m	F�vU��&�l	��$r� �� ���� tC�� tn��!ti��uf�F�.��uf�F�#��uf�F���uf�F$����&�>:	� f����"u&�>m	�t� � &�>m	�w�&�>m	�u%���f  � ���"tf��#ta�� u&�>m	�t
&�>m	 t�f%�����uf�F�9��uf�F�.��uf�F�#�� uf�F���uf�F$����&�>�	� f��]fX�N�]�n�^fXf^f[f`�^�  �(���&�  t�2F�v��&� F��&� F�� �
������������������������@BDFH�L�����������dF���3s� .��%
���t&�  .����e�� &�& �&	 F�G�� ��&�  t��� �ڻ  �ջ@ �л� ��F�v� �ۋ^���� �^���>� �� &�  ��ul��� �^t��l�>�F�v� �ۋ^���� �^���>� �� &�  ��um��� �^t��m��F�v^V� �ۋ^ ���� �^ ���>� �� ��&�  un��� �^t��n���F�v^V� �ۋ^ ���� �^ ���>� �� ��&�  uo��� �^t��o���܃��t"6�?�t&�  f^f[f]��fU��&�6 �&�  tA� �F t��6�76���t&�  tA��*�             ~��ۇۇۇۇ�fUj �jfUj�dfUj�^fUj�XfUj�RfUj�LfUj�FfUj �*fUj�$fUj�fUj�fUj�fUj�fUj�fUj� ��fSf�   ��ۇۇۇۇ�f��fSf3�fV�� �޾  f��f��g���  ^ ���F �� gf���  ����,��,fPfRf�^(f�F,f�^�f�F f�^ f�F$f��f�F��^�����f����f�^,f�F(gf��H	  gf���  ��(6f�W$f�V$6f�W f�V 6f�Wf�V6f�Wf�V6f�Wf�V6f�Wf�V6f�Wf�V��f��f�V�  f�Vgf��    fBg��    g��P"   gf���  g���  (fZfX��gf��H	  g��m   �� gf���     �� f�^���^Pf�vf���Fg�CC�Fg�CC�Fg�%���FXf�^��� �# �� .g�]  �^�  f��g���  �^�gf��    �^f���^f^f[��f]fϻP ���H�� ���]�f�^���^Pf�vf���=g�CC�  g�CC�Fg�CC�O��fSfV���� �۾  f��f�����fPf�F�f�Ff�F�f�Ff�F�f�FfX��������f��j j h�fUf��PfSfV�� �  ��f��f����Çۇ�fU��j!h� �e�6��t e�6�� e�6�
� e�6��Y�� ��H�N�� ��ef�>T	����f��g��*  g��,  g��2  g��4  f  ef�>H	f���)  gf���Q��f]f�fU��j%���fU��j&���fU��j*���fUf��=Jtj/����rf]f�fU��j3���fU��j\���ۇۇۇ�fPfS�� �ظ  f��f��gf��H	  gf��    gf��X"   Kg��    ��(gf���  f[fX��f]��$��fχۇۇۇۇ�fUjP�(fUjQ�"fUjR�fUjS�fUjT�fUjU�
fUjV�fUjW��fSfV�� �޾  f��f�����/��ۇېfUjf��fSfV�� �޾  f��f��gf��H	  gƃL  g���  ^ �����   f`��P �ػ�ù� ��� ��f3� �"�f��f��&g��     ukf�0gf�]6  gf�<]2  �60�t&gf��        g�]6   ہ� �f߃�g&gf��    f��g f�   �f�f   ����xdgf�f�:f�>&gf��    �� �f��f��
f��gf��f�Bdg�  �J dg��^�F�N �f��ef�X	f�Pdgf�Sf�Hf�Tdgf�Sf�L� �"��fa����fPfSfR��P �ػ� ��� ��f3�f�Bf�tNdg� ��f���F�� 	^f�>f�:dgf�ef�X	f�Hdgf�Sf�Ldgf�S �"��F u��fZf[fX�fRf��   sLgf�f��   v>fPfS �% �&gf� % �gf�f��f��
f��f��
f��+�B&g�� tCJu�f[fXfZ�f��f+�vf����f��   f�f�f+�w�f3���fP� ef�>� t�  f����dgf��� fX�e��@ � �fPfQf��   dgf������gf��X  ��fYfX�fPfQf��   gf��X  dgf��������fYfX�V3��V� � �u���Ƅ� �^À����t���^�u�ø �  �(V�6`�V�6���Q�t�ȃ�������u���
�D u���Y^�V�6`�V�6���t#Q�ȃ�������u��������Y^��^�V�6`�V�6��q�tDQ�ȃ������Y�L�d��P$�<�Xu�L � t�L �u�d��t�L�t�L@�^�V�6`�V�6���t#QP� �u�=�M�����������XY^��^�V3��V� ���tƄ� �^��^�PV���3��
PV���� �t
Ƅ� Ƅ� �^X�V�6`�V�6���tQ� ������Y�^�VW3��6`�� VW3��6p� VW3��6�� VW3��6�� VW� �6�� VW� �6�� VW� �6�� VW3��6`� VW3��6p� VW3��6�� VW3��6�� VW� �6��yVW� �6��nVW� �6��cV�6`� V�6p� V�6��~V�6��wV�6��pV�6��iV�6��bfPfQR� �������t�d���D � �L �z���ufPfQR�z �������t�d���D
  �@�L �H��CWfPfQR�G �t�d���D �D�L � �D t�D�f�Lg��~  �*DD���ZfYfX_^���PQV���6`� � ����6�� � ^YXèt�� �������f`�ts�&l��l tf�|��  uf��f�D�&l���D uIg�FfQ�D  tf+��fYref��   t'f��f�f��   v�D u�D@ uAf;dw&�� �D  tf�����L�L���mfa�f��
������ٸ �(� �  �(PQ�L����� m�t s
�ts�� YX�PR�D tef��   t3��D� � ��1 �ZX�PR�D tef��   t3��D� � �� $��ZX�S�\��n��$[�fQfRfVfW�l t�l t�`��������l�L�D t�] �D  tf+�f��f�>h��f�hf_f^fZfY�fPfQfRfVfW�D t�% �D  tf+�f�6hf����&l�f_f^fZfYfX�f�f�LfAf�   �D u*�|rf�   f��f����f��f;�u	f��    �f3��D� t�f��ef��   t����D u�|r
f��P3�f��Xf�D��D� t�ef��   t���P�d��ef��   uZfSR3��� f�\����D�D���~�D�����D�D	�| u�D tg�]�  �D�g�]�  �D
�Zf[X��D t��D �� � �D�� � �D�� � �D�� � �D@�� � �D�� � �D	�� � X�SR�D t�@��> �\����Z[�SR�D t� �"�" S�\����[�t�T���*T����Z[�RW�|��v�
�t����_Z�PfQfVfW�� �����g�#�� tg&�g�f���� tg&�g�f���gf&�g�f_f^fYX�fSfVfW�� ��f��f��� fKfPf��f��f��f;0s&g��     t
&gf�4�    �� �fVf��   f@f;�w.f��f��f;0s&g��     t
&gf�<�    �� �f;�t�fXf[����fNf�t"f;�r9f��uf��t�f��uf��fJf�fB�f3�fFf+�f;�sf�����f_f^f[���fPfRW����� ��&�{ �P ���� ��>`2�ef��   t������ � f���� � � � � ��� ���f�f�f3�ef��   t��f��� � �� � �����f��>p2�ef��   t������ � f���� � �� � ������f�f�f3�ef��   t��f��� � �� � �����f��>�2�ef��   t������ � f���� � �� � ������f�f�f3�ef��   t��f��� � �� � �����f��>�2�ef��   t������ � f���� � �� � ������f�f�f3�ef��   t��f��� � �� � �����f��>�2�ef��   t������ � f����� � ��� � ���Ć��f�f�f3�ef��   t���f��� � ��� � ���Ɔ�f��>�2�ef��   t������ � f����� � ��� � ���Ȇ��f�f�f3�ef��   t���f��� � ��� � ���ʆ�f��>�2�ef��   t������ � f����� � ��� � ���̆��f�f�f3�ef��   t���f��� � ��� � ���Ά�f�2���� � � ���� ef��   tZ�>�&�M f3��4�� � �� � ���� � ��f��3��� � f��f��f�f�f3��T�� � �� � ���� � ��f���_fZfX�fUf��jPh� �h0��&l�e�� u��u�lj��
��� f����  �&��������&�?�6����&��f�Nf��f�f�d� f�>� tf��df�f��    f����r��f3�f��s	f����C������g�]$  ��t �$����d�6�Ĉ&2���� �6�&2� �� ��&��	�&d��&$f���ff�
��d*�� �&$f���f��fPf;dvf�
f�   ��wf��f;�w�k�re�&���f;dsf�dfX��f��f���6$d �&�f�
f���^f���
�6��f]f�f]f�VQ�6`� �D � ������Y^�           <tCf`f��gf�e�h� <r�f%�   g�EJ  gf�]�6g�Cg�e�
�tg�Mfað�����u%�� �>d�6f� � 3��l t� g�e�ðg�M�����t�� f���&g�C
  �f��f��f3�f��0   tf�   f��   tf���0�sX&gf�f��   t�f�tK��Gf;dv��<�.l s��0&gf�f��f��   t�Qf�>h���(&g�C
f�h&gf�C2������t��Vf���f�>h&gf9{t�� u&g�{
 t2�
�0&g�C
��t�
�"�l u���� t	��f���4��&l�2�����?�t�3��� f���&gf�{�&gf�3&gf�    &g�C  f��@   u:f��f3�f3�fQfP��f;�s&gf�D�&gf�L�&gffFfXf�gf)$fYu��w�� ��f3�f�f�f�tfIfPf��f��f;�s/f��f��f;0s
dgf��    �� ���&gf�T�&gf�   f@fFf;�v�fXf%�  gf�U�6g�Bf�t&gf)fY&g�s�	f;�w2�&gf�����?�u2�ð�����t��If���l t��9�f�d&gf;s��&�l�m&g�C
f�>h&gf�{�� t�r���2������t��4f���Mf�>h&g�C
�;u�l t�� t	�;f�����&l�2�ð
�����t��6f��f����f���f�>hf�&g�C
�� u&gff9dr�� �E�2�ð
ð�����t��9f��f����f��� f�>hf�&g�C
� u&gff9dr� f�����2�ð
ð�����t��%��s)��Br2���Bu��3��������l�ƇB��ð�����t��*��s.g�e���Brug�M@��3��������l�2��ƇB �ðá@@u@�@�;@�gf�]f��f��&gf�sf��&gfs&gf��fUf��f��jPh� �e�6�s�w�f��f]f�f��jK�F�      V�6`�V�6�Q�<��t�ȃ�������_��Y^�V�6`�V�6�Q���t�ȃ�������d��u	�t�L� �Y^�V�6`�[V�6p�TV�6��MV�6��FV�6��?V�6��8V�6��1V�6`�fV�6p�_V�6��XV�6��QV�6��JV�6��CV�6��<WfPfQR���t%� �L �D
�_��D t�D
�R�f�Lg�M�  ��A�WfPfQR�E��t�L �D�&��D t�D��f�Lg�M�  �*DD��      � F(�&q(�(�(")~)�(�(�)�)�&�&�)�&�&fPWfS3����ef��   t-�t)��f��<r� ��f���   f��g.���&  �f[_fX��f[_fX�fPfVfSfRfWfUf����ef��   �f�6`�ugf���   g���   g�E�� g���   �� gf���   f���   f�� �� f��@tcf��pt)f���   � f�� �� �gf���   �� �� �g�d>g��t�ug�L>�g�L>�@tg�L>� g�L7 �n�Ygf���   gf�<>g�Dg���   g�O �#�3gf���   gf�<>g�g���   g�O fCg:��   rf3�g���   � �f]f_fZf[f^fX��f]f_fZf[f^fX�fVf�6`g���   gƆ�    gƆ�   gƆ�   �f^�fVf�6`g���   gƆ�    gƆ�   gƆ�   f^�fVf�6`g���   gƆ�    gƆ�   gƆ�   f^�fVf�6`g���   gƆ�    gƆ�   gƆ�   �f^�fVfPfWfQf�6`f��� ��f��gf�<>gf�f�   �%fYf_fXf^�fVfWfQfPf�6`f��� ��f��gf�<>g�G tgf�Gf�   �� fXfYf_f^�fXfP�� � f3��� � ���� � ����fVfPfWfQf�6`2����f�   � fYf_fXf^�$<�$�r�8���,��$<�$�r�%�����fVfPf�6`f3�g���   g���   g���   g���   g���   g���   g���   g���   gf���   ��Z��\�fXf^�fPgf���   $� ��f��fX�gƆ�    gƆ�    g���   gf���   �  g"r-}8�p�����v--------�&-�&---------------------------------------------------------------------�.---f/----------------------------����4�4-�-���-----�-�---�-���----------------------------------------C-�-O-�-[-�-u-�-�-#-�-�-�-}---------------------------------
P%�W%w%�~%�%�%�%�%��%��%��%��%��%��%��%��%�&�&R�jPh� ��� s����.��`*���Z�ef��   t2fQf�   .g;�\,  t	��fY��P�����g.��^,  ��fY�ZÇ�P[���Z�tef��   �����        Y-.��wgf�e�fSf��g.�]0-  f[sgf�M���� �� �� f`jPfWfVfQ� f�p  �| t����fYf^f_��dfY�L�f���Tf_�|gf�]f��fXH�D�D�\
�\f���\�\�D��D�� h@3ۋ|&�;r;Dw������g�t$faË|+L���&��~�����D  �����f`jPf����=pr/-p=x s'3ɇL�" h@3ۋ|&�= r�9�����fa�����6 fPfWfVj�f���8$�f��f�f�f�f�f^f_fX�fQfWfVjPf�p  � �| t>;r:;Tw5;6 t��h@�L�|&9t�����f��f��h�.h8&�u˃���f^f_fY��u/ef��  @ u�À>N�u��>Lt�M�O��L �`�M�B��>N��N t��PSh� �&�ߨt�� ���`ef��  @ u3۸` �&[X��PS�t=�N<�uVh� ��vd�<�^u&�d�ef��  @ t<�u�L�3�<�u�` �� [X���u�h� $���  t�âPh� �&�ߨt�� �5�X��PSef��   u82�ef��  u���N ef��  @ t�` �Y �d �S 䒢�� �H [X�             PSV��  ���:h�� �E ��h ���� �7 ��h ���|��^[X�� �PS� ��h ��[X�PS� �Ё�h  ��[X�Q�ȃ����ظ ��Y�    fU��f��fR�� �ں  f��f����Otv���t-gf���     t���w���r	2��N�H�fZ����j��g���  rf���Zf;T u�f��f���F tgf���  @   u��~ �fZ��f]f�<R� <Su�fR�@ f��f��Sg��   ����[fZu�<R�& fSf�^
f��f^�f[�i�gf���     �Z�gf���     �J�f�~
 �  �>���fPfSfQfVfWf���F  �F �� ��Á� ��rf�^f��f��fދ���Hg9C�Ug9C�Mgf�s�s�N�� �N gf�s�qs�N�� �N gf��T	  gf�sgf�{gf���   gf���   gf�sgf�{gf���   gf���   ��  ��� ��  ��� f����f��g�sf����f��g�{�F�� �vs:g���    u�Ng�� 	  t�N�Ftg���   g�� 	  ��N �+f����f����� tg�g����gf�g��F t�Ftg���  ��Ftg�� 	  ��f_f^fYf[fX�f �N@�f�
�t�f��N��F �SR����x���Ft����` �Fu��wglB�����{wgnB���K �Z[�t�gf���      tg�~�u	g�~�u����g�~sg�~v	g�~ u����P�a�F �aX�P3��F �aX�f]NNg�g��a��䀆��a��䀆�$��a�F �����fWfVfPfQg���   �S gf���  f��f��g�?Mtg�?Zu7f��gf�Of��f��f�g�
tf;�� f;�� f��g�?Ztf����fYfXf^f_� 6�t�W�U�������tH�V慀>U�u5< u	�>Wu*�1<u$�>W w3ۊW���u.���4r�f���N�U������뺀 ��ef���   t�Sރ�Z[f^f[f`�^�        P���P �ظ� �踀 ������U �V��W��9�� �� ����X�P��� �ظ0���� tNd�1 ��8 ��&�>  �u&�  �&�>~  �u&�~  �&�> �u&� �&�>� �u&�� ��X�� �* �fSV�� ��ƃ��df�\f��d�\f��f��^f[�fS��� ��fPf��dgf��    f�� ���fXf%�  f��f[�� �fPfQfW��� �ظ� ��f�   �� 	uf3���  tf��f�   � &gf�$�    �  &gf	�    Gf   Iu� �"�f_fYfX�h� �&{�� �P��� �ظ0���� tV��@ uNd�1 ��8 ��&�>  �u&�  �&�>~  �u&�~  �&�> �u&� �&�>� �u&�� ��X��               �7�7�7�7p8@9 ::�: ;0;@;P;p;�;�A@C�C�D�D�E`FG�H�KL�L�L�N�N�ۇ�f`�����^s���@re�>	t�.��7fa�=��t�F����F������F�F�e�6 �F�F  �Ӈ��F Çۇۇۇۇې�?'���^�F e�>��t��F�Çۇ�e��- ���F�s�F�F Çۇۇۇ��tWe��- ��;�rO�-rT��3ҋ:f�6�(� B��<�t�B;�r���F���  �D  �R��Zre���V�F ��F����F�������F���ۇۇۇۇۇۇې�F �>8�� f��;>='�� ;:�� f��f����f�(�?��� �f��?'����f>$���t1���us��;Osk��f�7���f6 � �gf&�g�� �"�Çۺ f��g gf�g�f�gf�g�f�gf�g�f�gf�g� �"��,�w�<w�R��F����F����F����ې�F ;:�� f��f�Ӹ��8��(�� ��f�(���=���s e���u�e��f3�f�>�(gf��gf�L�f��3ɇO�>�e;�ue�>���f> ��e)������3�&gf�'sA&g!f��Kt�������Ý�F����F���ۇۇۇۇۇۇې� �@�FÇۇۇۇ��F e�>��tR;:sRf��f�>�(g�<��tB� ���(���u=f����f>�(ef>H	f�6?'��f6$� � gf&�g��Iu���F����F����F����F e�>���s ;:ssf��f�>�(g�<��tc�����(���t^f����f6�(ef6H	f�>?'��f>$� � gf&�g�gf�g�f�gf�g�f�gf�g�f�gf�g�Iu� �"���F����F����F���ۇۇۇۇۇې�F�Çۇۇۇۇې�F�Çۇۇۇۇېe���^�F Çې�-rf��f��(g�\����^�F Ç�f�F&f��f��f���e���Nf3�Nf��(Fg�<��t�&g�7f��g�D���&g�f���ޝ�F Çۇې <3< <�;�ۇۇۇ�<ss�F f���.���;�ۇۇۇۇۇې�@�FÇۇۇۇېf�F&f��f��f���ۇۇۇۇۇېf�F&f��f��f��}f�vf�F$f��f���F��   �<�<`=u=�=�>?<?J?�?@-@<wr�(���f`f��f��g.�EP<  fa�ef�	g�Eg�E �gf�}&f��gf�E f��B�� ��f3�f�   �gf�f%����gf�g���ef���˃�g gf�g�f   ��gf�E&f��f+�g�} gf�}$f��gf�Ef�jf�(  gf�g�gf�g�f��   gf�g�gf�g�f�  gf�g�gf�g�&g�G�&g�G�  f��  gf�Eg�E �f�,f% ���gf�Eg�E ���f��f��ef��e+�e+�f�gf�Eg�E ø��e��e+�e+��  ef�6�ef�>�&g�,�����
smN;�u�ef�6�e;6�vv� ef�>�e)�e)�;��5 ���f��gf�4�����gf�<������gf&�g�� f3�gf�~��gf�g�f��&g������ e��&gf�������� ��F f�V�e��- ��e+�� �� ������|����V��� ��� �����B��F��ef�6�ef�>�;�tY����� ���g&gf������%��f;�tN;�u��3N&g�$�    ����ؚ
(e���F f��s�P �ظ� �����F����� s%�� ��f��&gf��    f�� ���gf�Ug�E �g�E�� �gf�Eg�E ø� ��gf�}&f��gf�E f��!�&gf�f��!�&gf�f��!�&gf�f��!�&gf�f��f3�&gf�f��&gf�f��!�&gf�f��!�&gf�f��g�E ø� ��gf�u&f��gf�E f��gf&�#�gf&�#�gf&�#�gf&�#�gf&�gf&�gf&�#�gf&�#�g�E �e��g�Ee��g�Eg�E ø ����e�>�t2e�>�Pt*ef�6�� &gf��        &gf��       fF��e������ ��P�� � f��&g��   H &g��   �fF��f��&g��     F&g��    �F&g��    &F&g��    ,F&g��    2F&g��    8F&g��    >F&g��    De�>�pt2e�>�Pt*ef�6�� &gf��        &gf��       fF��e����p�� ��P�� � f��&g��   H &g��   �fF��f��&g��    JF&g��    PF&g��    VF&g��    \F&g��    bF&g��    hF&g��    nF&g��    tg�E �      0B�BB�ۇۇۇۇ��F <s(���.���A�ۇۇۇۇۇۇ�;='w�����^��F����F���ۇ�f�F&f��f��f�f�v$f��f�Ff��f��g&�gf�g����7;='w2f�$f3�g&�
�u)��g���'  �t&gf��2�f�gf�g�f3�Iu���F����F���ۇۇۇ�f�v$f��f�Ff�gf&���f��=�uY�V;='wQ� f��f�$U�g gf&�f�����'�t92��&gf��Gf�&gf��Gf�&gf��Gf�&gf��Iu�] �"���F���]�F���ۇۇۇۇ��F <s-;:s-f����f�(g�:�tf�v$f��f�^f��<��F����F���ۇۇۇۇۇۇې�F ;:� f��f����f6�(�<��� ����� �L��+�|b�� �����\e)�f�<�e;>�u+�|e�>��+�|��f> f�   3۸��&g�&g!����
�f�Iu�
�te��`e��- ��;�rSe��- ��e+���;�s	��+��Lr<����f�<�\�e;>�s+�f� ��e�>��<�e�>����
r���F����F��\���^���F���ۇۇۇۇۇۇ�<wr
�F �F �
�F���F�Çۇې<r�F�� ��� f��< t^f��f�v$f��f�Ff�gf&�f��gf&�f�6�(f�uf�t�:f3�gf;�ugf;D�tB��gf��gf�D��F �@�F��:f�F&f��f��f�h� f��(gf��&gf�f��gf�D�&gf�f���F Çۇۇۇۇۇۇ�<wr�:�F�F � �F�� <taf�F&f��f��f�h� �:f3�f�6�(f��(g�<��t%&g�f��gf��&gf�f��gf�D�&gf�f��C��e���F�F �Kf�v$f��f�Ff�h� gf&�f��gf&��:f3�f�>�(gf;�ugf;D�t	B���F���V�F Çۇې�F <sr;:srf����f�(g�:�t`f�~$f��f�^f�&g�w&g�7&gf�wf��&gf�Of�&g�OfW��f_YXr:e�� tU�nf��f�N�F]��F���F��Pf3�f���pX&g�&g�GÐ0G�G�G`G�ۇۇۇۇۇ��F ��<s
���.���F�F��C�F��=� �*&g�?�u�&g�  u��F  � �f���
�@���@ �F�F �&@��Çۇۇۇۇ�;:s�f����f�(g�:�t�f�v$f��f�Ff�&g�v&g�6&g�~	 tD+&@f��ef>L	fV��	f^f��&gf�wf��&gf�G
f�&g�O	fRfW�
f_fZ�s�f���@���Z
fV�	f^&g�~	 tf��f��ef6L	fW��	f^&@f��&gf�wf��&gf�Gf�&g�OfW�a
f^s	�@�
�������	&g�G&g�Gf�   @&g�;&g�&g�D;&g�G&g�D;&g�G&g�D;
&g�G
&g�G�&g�G  Ð<r�F��gf�^$f��f�Ff�h� &gf�f��   v�F��>f�u�F �3f���; r*f��f���/ rf���� �~ t< t�F���$��o�LÇۇۇۇۇېfRfVfW&g�;t8r�F��� &gf�Cf��&gf�Sf�f�f=   wf+��� �F���{&g�S�rqf��&gf�C���u��f�>�(g;D�r�F���K&g�S�� @r�F���9f�f���  f���g;D�v�F���+�g�- f��&gf�Sf���f_f^fZÇۇۇۇېf;�w� f�f;�wf+� �f+���f�f;�wf+�� �f+��Çۇۇۇۇۇۋك�f��g�&gf�&gf�&gf�f��f��fIu���&g�&g�&g�fGfF���F Çۇۇۇۇۇۇ�<t�F �+�F��� t� �f�fOf�fNf��f��f�� tf��f���ك�f���gf&�g���= uf��f���g&�g��Çۇ�fRQWf�Ѓ>F uH��ǋ>D���B������>F&f�= u��t�����Bf� f 0  f��gf�f   ��f�F�D�BI��+�f��f�_YfZÇۇۇۇېfPQW3��>F�t ����BI��+�����Bf3�f����_YfXÇۇۇۇۇې�F <�; w@f�F&f��f��f����� �<+���f���':�tf����gf�g���Iu�='�F��F����ۇۇۇۇۇۇ��&` r�F��c<tr�F��W���Rf�F&f��f��f�h� � &g�f���XH&g�f���@&g�f���  &g�f���  &g�f���F Çۇۇۇۇۇۇ�<wD�� w:f�   �:f�>�(g�<��t	F���F��$g��  g�D�  �ve���F �	����F�Çې@M�MM NpNMM%M%M�F �&` s3<	s5���.���L�@�F��F ��� t�F���� t�F�� ��F����F���ې�>�( u&f�4�F f��f���^6�Gf��f�f�� t�C��(�FÇۇۇۇۇۇ�:Xsz������p+ut
�u~f�F&�6f��f�v �64f�f�ta&gf�@uRf��=�uIf�@+�f��ef>L	f�׊����gf&�g��̀���g&�g��f����&@��F����F����F����Çۇۇېf�X3۰��p+< t��Iu��F��/e�>��� ��r+f��t+f�6 &gf�6�� � �gf&�g����^Çۀ� t:�(t!:Xs2���� ��p+< t��F��>Xt��F����F Ë�f����<wctB�.`rh� &f�lf�\�Vf���V�f;\u1�F <t�.` �+�6` �#f;\u�6`�.` �F �
�F���F��     ��e��- ��e+�;�rWef�>�e��+���+�r8\�<�t�<e���e��<�\��� f� � &g	��Ku���Ý�����j 딝S+�� [s��� �e��e+���;�r�r���� �Se��- ��e+���e��e+�;�v� �[Çۇۇۇۇۇۇې� �SV� � f� ��ef�>�� &g�T��u+�;�r��e���+�+�v3;�s/� &g�T��t+�;�r����W&g�T��u+�;�r�[+��	 �+�w�^[ÐfPfQfRfVfW��� �e;>��� +�Sf�6(f��� &gf��gf�g��+�u�[V����f�ef��+�e���+�f����f+�f���gf&�g�f�6(f�   ����gf&�g�gf�g�%��f�gf�g�f�gf�g�f�gf�g�Iu�^f�:f��(g�L�����t;�r+�g�L��Hu�f_f^fZfYfX�e��- ��e+�+�s	��S���[�� �e��- ��e+�e��e+�v��P��� ��[�Ð;:sf��fPf��(g�<��fXt���F��Çۇۇۇۇۇۇې��f��Hgf�g�f�$f�='gf�4M='  gf�4�gf&�g�Iu�Çۇۇۇۇۇۇېgf&�@uUf��=�uL� f��f�='gf�<M='  ��f>$gf&�g�gf�g�f�gf�g�f�gf�g�f�gf�g�Iu� �"���F��Çۇۇۇۇۇۇ�fP���wU�nf�~f��Ff�Ff�]fX�je�e�>����f�E�Ef��ef�>�f��Շۇ��r;='�� gf&�f��f��f���Fta
�uv�����'�tl����f>$���tt���u_��g;ZsVf�f�ޱ��g2��f6 �gf&�g��f���Iu� �"��Çۇۇۇۇۃ>8�[ ;>='� ���?'���F��=��F��6�ۇۇۇې� f��g gf�g�f�gf�g�f�gf�g�f�gf�g�I�.�� �"�Á�� w��� ��v�뤇ۇۇۇۇې����f��t+f�$f��f��
f�f��  @ sf+�fǜ���g&gf�8f� &gf�8��(e��%  9�r+u �"؝É�r+f�   �e� 	uf3�e��  tef���� �g f�   f�   � &gf��f�CIu��    SQRfV3���f�6�)f�t&gF;�s&gf�6��+؋и �S�;�s�����f^ZY[�f`��3���f�6�)f��� &gF&gf�6f�u�^;��� e��e+���;��� f�6�)f� ef�>�gf�<�&g�N�d;�v��+�&g)NS&gf�^��g&gf�V�f��f��f�gf�g�f   gf�g�f   gf�g�f   gf�g�&gf�TV��&g�V[�t
&gf�6뎝�f+> ��e�>������^+��C���=�fa�f`f3�f� ��ef�6�e��;�vK&gf�d��s�����t2;�v3&gf�d��r���� &gf�D��&gf�D��&gf�D��NO��붍|��ɝ�����ef�6�e��;�v&gf�d��s����e��e�6�gf�<���+��� ��f�6�)&gf�^�&gf�f+�r@f��&g;F
s5��&g�V&g�TF&g�Ff3�gf�g�gf�g�gf�g�gf�g����<f����4f��&gf�&gf�6f�uf�6�)&gf�^f;�t�f+�r�f��&g;F
s�뗝�fa�fVfW��sf��)��� � g�]�)  e��e+���;�s�ع f��@gf�E   - r���
���ٸ������ f����Agf�M   f��gf���  �� �f��f��
gf�8f+�f��&gf�    &g�W&g�O
&g�O&gf�_3�fWf���g�g�@�����g�g�f_����)f�6�)f�uf�>�)�f��&gf�6f�u�&gf�;����f_f^�fSfRfV��ef�H	f�ð)  f�6�)f�t2&g�F&g;F
u&gf�&gf���)�&g�V��ֶ�f��&gf�6�ɝf^fZf[� 6X�X�XfPf���P �ظ� ��f��g.�EX  fX�fSfV� dg�C��� �1�dg�{rdg�C����^�f��dgsf^f[���� ��� ��fS�P ��f[�fP�F�u<�u8e�>`	e�b	��
s�� r e�b	 ef��   �&�  �v��	fXù����fPfQf� f�   gf�M   �t
dgf�    ��f��   fYfX�fPQdg�  e�b	dg�Cf�\dgf�C� �XI��p+udg��:����dg�{r,dg�e�>� � dg�ef�>�   t�>c+udg�YfX�fUfPfQfRfW�� �¡@dg���  dgƃ�   f3�f3�f3�dg�D;
 dg�D;�dg�D;��dg�D;�dg�D; �f���t�2�dg�{re�>� r�f���� s�f_fZfYfXf]�fPfRfWfUQfV���dgƄ3�   dg�{�
 e�>	��� f�>�(f�.�(�:f3�g�<���� fXdg���  fPdg��3�  dgƄ3�   dgfǄ3�      dgfǄ3�      g�D���dg��3�  gf��f����dgf��3�  >gf�D� f�u>gf�D�f�t,>gf�D� dgf��3�  >gf�D�dgf��3�  dg��3�  g���(   udg��3�  dg�f��BI�,���Yf]f_fZfX�fPfQfRfW�  f����dgf��3�  dgfǄ3�      ef��f=   tf�$f   �w�dgf��3�  dgƄ3�   f��f3�� �f���t%dg���  dgf��3�  dgf��3�  ��f���f_fZfYfX�dgƄ3�   �fPfQfWRf��dgƄ�   ef�>��tWf��dg�?Mtdg�?ZuEf��f��@dg�Wdg� udg���  dg��3�  dg��3�  ��dg�?Zt�f��f���Zf_fYfX�fVfWfQf��gf���  �f�6d	�� g�g�fYf_f^�fSfVfWPQR�� ��f��f3��@ dg�D7
t)e�>	�u!dg�D7dg�\7dg�T7f`����fa
�uf�����ZYXf_f^f[À��t����fRf�����dg�{re�>	�u��f��gf���'  fZÐfRfVfSdg�D;dg�D;
�� �v<sdg�L;
f����&gf��    f����Ƌ:If����f6�(f�Tf�4���t%��f���tJ��&gf����f��f;�t�u��u�����f[dg�L;dg�T;f^fZ�fPfQRdgfǄ3�      dgfǄ3�      dgfǄ3�      dgfǄ3�      f3����� ��dgD;���� t<&gf��    f��	s�] �&f��f;�t�O P� ����dgD;
Xdgf��3�  ��BA��r���dg�D;
�tdg���  dg�D;dg���  ��ZfYfX���P� ����dg D;� ��dgD;��X�fSfRVf� e;>�s?dgf����� u�f�   f��f�� @  e;>�sdgf;�u������f��^fZf[�f�������fP�U f�>�) tJ� �Y�fWef�>�
f��f���  �Ff����dgf�Ge��
f���Bdgf�Gf���F��f_fX�fPfSfVfWQf�6$ef�>H	f���)  f��   �` dgf��f��f;�uC���%f��)f;�� f3�dgf�f��Cdgf��f����e�>�	Yf_f^f[fX�fPfRfWe�>� �� ef�>���� f��dg�?Mtdg�?Zupf��f��dgf�W��dg� uDfPfRf��f��f�f�  f��f��f+�)f+�)f;�sgf���)      f@f;�r�fZfXdg�?Zt�Hf��f���f_fZfX�fPfVQe�>	t9e�>	t1f3��='gf�u?'  f+�)rQ� gf���)      f@��YF��Yf^fX�fPQf��   f+�)gf���)      e�� �- e�>� v$e����f��   f+�)gf���)      f@��YfX�       1a2aTa.cQctc�c�c1a1a1a1a1a1a1a1aja>bjPg.�M a  �À>c+u;d+r�c+ � ó�3�����3���>c+t	�c+� ó�3������ ��3�ef��f��dg�9Mt	dg�9Z�� dg�y udg9Yv	dg�Y;�sdg�9Z�~ dg�A@f���rpf���f����f��@Pdg�Adg�Qdgf�AUMB dgf�A    +�v6K�Mdg�f��A�f��dg�dg�A  dg�Ydgf�A    dgf�A    � [��ӻ� �t�� 3������ ��f��If��dg9Q�B dgf�yUMB �4 dgf�y    �& dg�A  dgf�A    dgf�A    � � 3���3��� ��fPfSfQef��f��dg�8Ztodg�8Muhdg�x uJdgf�XCf��f�f�dg�x u1f�dg�dg�dg�KAdgHf3�dgf�dgf�Kdgf�Kdgf�K�dgf�HAf��f�dg�8Zu�fYf[fXÃ>`+� �: �� �`+ � 2�ó�3�Ã>`+ � �D �� �`+  � 2�ó�3�À>b+� e��  �	 e�� ��e��
� 2�ó�3�À>b+ �5 e�>�
 �1 �3 e�>�
�
 �� 3����	 e�&���=�e��
� 2�ó�3��3�e��  � � 2��   �b�!�ÿ� �g� L�!    .� �      EMMXXXX0 WVSQR3��ء��t'���  �ؿ ��� �% ��u&� @.� .� ZY[^_�� =�# �!rI�ظ D�!r@� t:�D�  �!r0<�u,�D� � �!r= u�> %u�! ��� �>�!� 똴>�!����g=Z�� u����.�>`s�VPSQR� �	�!�� 2���ڴ�u2��;�t��t��2����u�ZY[X^�  Press any key when ready...
$EMM386 not installed - incorrect DOS version.

$
MICROSOFT Expanded Memory Manager 386  Version 4.49
Copyright Microsoft Corporation 1986, 1994

$  Available expanded memory . . . . . . . .       KB

$Expanded memory services unavailable. 

$  LIM/EMS version . . . . . . . . . . . . .   0.0
  Total expanded memory pages . . . . . . .     0
  Available expanded memory pages . . . . .     0
  Total handles . . . . . . . . . . . . . .     0
  Active handles  . . . . . . . . . . . . .     0
  Page frame segment  . . . . . . . . . . .  NONE  

$  Total upper memory available  . . . . . .       KB
  Largest Upper Memory Block available  . .       KB
  Upper memory starting address . . . . . .        

$EMM386 successfully installed.

$EMM386 Active.

$EMM386 Inactive.

$EMM386 Inactive.
Expanded memory data is inaccessible until EMM386 is re-activated.

$EMM386 is in Auto mode.
$Weitek Coprocessor support is enabled.
$Weitek Coprocessor support is disabled.
$Weitek Coprocessor is inaccessible until EMM386 is re-activated.

$Invalid parameter specified.
$[HMAon] is an invalid parameter on this machine.

$Insufficient memory for UMBs or virtual HMA.

$Page Frame Base Address adjusted.
$Mapping Register Address adjusted.
$Size of expanded memory pool adjusted.
$WARNING: Option ROM or RAM detected within page frame.

$WARNING: EMM386 installed without a LIM 3.2 compatible Page Frame

$WARNING: User specified ranges overlap.

$WARNING: Weitek Coprocessor not installed.

$EMM386 not installed - insufficient memory.

$EMM386 not installed - incorrect DOS version.

$EMM386 not installed - incorrect machine type.

$WARNING: Unable to set page frame base address--EMS unavailable.

$EMM386 already installed.

$EMM386 not installed - XMS manager not present.

$WARNING: This version of HIMEM.SYS may cause conflicts with EMM386.

$EMM386 not installed - other expanded memory manager detected.

$WARNING: E000 page frame address not recommended.

$EMM386 driver not installed.
$EMM386 Active.
$EMM386 Inactive.
$Expanded memory data is inaccessible until EMM386 is re-activated.
$EMM386 is in Auto mode.
$Unable to activate EMM386.
$Unable to de-activate EMM386 as UMBs are being provided 
and/or EMS is being used.
$Unable to place EMM386 in Auto mode.
$Weitek Coprocessor support is enabled.
$Weitek Coprocessor support is disabled.
$Unable to enable Weitek Coprocessor support
$Unable to disable Weitek Coprocessor support
$Weitek Coprocessor not installed.
$Weitek Coprocessor is inaccessible until EMM386 is re-activated.
$Turns on or off EMM386 expanded memory support.

EMM386 [ON | OFF | AUTO] [W=ON | W=OFF]

  ON | OFF | AUTO	Activates or suspends EMM386.EXE device driver,
                   	or places it in auto mode.
  W=ON | OFF		Turns on or off Weitek coprocessor support.
$Unable to turn EMM386 ON - protected mode software already running.

$Invalid parameter - $EMM386 not installed - protected mode software already running.

$EMM386 not installed - User requested abort.

$     �ʎںp�	�!�W�Ȏغ&�>	��� &��- &+���&+����� �� ���	�!�@2�����00�h�GG�ĈG&��- ��� ��� &��- &+���&+�� ��� &��� � �z &��� �3�m &�>��t&���f� � �EH�:�	�!&�>� t3�0������ �6 �)������ �' &���
�p �EH�q�	�!_� 
 d �'� �PSQRV��N��2��3�.��m��
�u�u� �0��G��݊�$0�G^ZY[X�0123456789ABCDEF� �PSQR��й �����.����G��}�ZY[X�               f`f3�f3��='�>8u� �� �@��( �p+fa�     H	Y	�	     onoffautow=onw=off/?;=@DHM                    PRW��w�>qt�su��
�u�)	�5�/�5�s� .� �������Ȏ�� �sth�>gu2.� ���� �Ȏ�� � � ���� � �%�s5��	�� �>iu�t����s��	� �>ku����s�>
� �st1� ���u�� �>mu����s��
�y���s��
�l2����2�= u�t�= rP��	�	�!X- ������0�	�!�>t t�l	�	�!� �r�t�e
�u��
�	�!�>t t�9�	�!_ZXú|�	�!����	�!&�&�E
&�E$+����	�!��SV�6� �m �t6�s�8 r/Ǉg ��w�su�s���w�su
�s�^[Às��W�ˎ�3�;�[u��OV�Q�Y^t
CC��u����_�VSP���3�&�G< t�<	t�O&�<t!<
t< t<	tGA;�w�<Ar<Zw �F��X[^�   �$�������������f���F �� �
�� ��!�h"��"��#�[$�=#�� �a$�#�$�$�                                               	
                                                                                                                                                                                                                                                                                                                                                                                          � �                                                                                                                                                   �? ��� ���                                                                                                                                                                                                                                                                                                                                                                                         � � � � � � � � � � � � � � � � � � � ��                                                                                                                                ON OFF AUTO FRAME=ROMCOMPRESSVERBOSE ����������                                                      SMARTAAR CACHCMPQ                                  ����                                   � �TOSHIBA  �� �03COMPAQ� �ZDS�� �auto�n>�9�kb6j�
����*.�\.�&^�1�Ѝ& SRUW�츭�؋^�Ë^
&�G  �  &�G&�G �	.�U�as�i�f��s�Z�  ��&��
s�S� ���&����Z藟���ظ  ��������sef��   �G���t#
�u�@�g�uef�� �  �'ef�������uef�� � �jj3����jj� ��3� e����3� �@f3��f�   te� 	�H�^�Ë^
&��r�����t.��ef��� ���3� ���r�t
ef��   ���ef��� �r.f�Af��
f��f��
f�f p  fd.f�.f��f�.�>�uf   �=f�f   ��8f�,f�  f��f�0f�u
ef�����9f��
$�f= �  v� �.;As.�A.�>>uef�� .;?s.�?.�>=uef�� ���ef��� t� �ʋef��� �� �eef��� �� �ef��� �y ���ef��� t�h��zfef��� �V f3���8e��
e�� e�&��e� 	te��e�	e��<u
e�>� t�<ue�
 $��   ��e���  ��f�>� u.�>�u	.����f�   ��f�   f��t.����ش	�!��f����f��� �cf�>� t�����'腔3����  f���Z&f�T f���  f���&f�d f���� ��f����&f�� df���� f����&f�,df��&���&��  ��M�����f3��P.�U? f��A Z;�s
ef��� ��^�Ë^
&�G .�U&�G.�>��� ��������ش	�!�  ����� 	t-��� 	u�����ش	�!�>	u�&���ش	�!�`�>�t#�>�u�����ش	�!�K�� t�8���ش	�!3�_]Z[.�\.�&^�f�������6���]� ��ۺ���>������ش	�!��`�������ǎ߿��ǿ<���
���.������e�>	�t"e� 	te�>	 te� 	�
ef��   e�>	�ue�	 .�>�u .�>�t.�>�te�>	te�>	ue�	e�	 �%&�?&;Av%&�>=t
&�A&�?�&�A&�>>uef�� �n"e�>��u3e�>	t=e�>	t5�>8uef�� @  �ef��e�	�M�.�> - t
ef��   �a�PW�< t�<	t�3�<t<
t< t<	tA<ar<zw$ߪ���2��_X�f`���؋����f��$gg�,��  f�|�HIGH� f�|SCAN� .�����f�<MAONt;�<=�r�>$ �i�t�b��\= �U=� �Nd�:e���$��H���<=u�A�/��)=? �"��
d�d+.��� ���u�1諏��0褏
�u�ef��   .�� ���<H�m�<Pt��f��$gg�,��  <P��e�>����������.�>�t
� �<��e���.�>>��N����t� ��=@ s�@ �= �w�t$��� �ef�� .�A.�>�T�<=u*�>% �<�G�5��/=� �(@d�X�%��%f�|�LTBOu�|OTue�� ���e�>	�������� ���e�	���>& ���<=��������!�����= ��;�v���% �f3ۻ  f����f��f���  f�� ���;�r��H.��@��d�<�&��tf�<MAXTud�l���_�>' �L�<=�Ef3��M�;��5= �.= �'f��
df�d�'�� e�>���N��� ���f�<NONE�;�e�	����f�>�����<=�������������u��������f�|�NOMOu%f�|VEXB���|DA��ef��   ��	�f�<OEMSue�	���zf�<OINTuef��@���df�<OPFC� .�����Mf�<OA20uf�|TRAPuef��   ���*f�<OVCPu�|Iu.�����f�<OHI � .������f�<OTR ��.�������<IN�L ���<=��.�>=�������� � ��= �� �t$��� �ef�� .�?.�=�e�>���y��r��l��f= �_����H��؁��e���Re�>	��>N�޿�� �u	e�	 �2��� ��e�	���
= v=� ��
���-� �؀������|�=���>�����.�>�t
� �e���� �����������f�<MSINu�|TSu��ef�&������f�|�EMS=�}�����*f�|�ROM=t/f�|�RAM=t�<OMt)�<AM�Q.�� ���N������ ������ N.���>�� ���!N�< ��<0��<Z�.�� �� �<=�7 e�>	��� F�޿�� �u	e�	�� ��� ��� e�	 �� f�|�WIN=�� ���&�\��<=�� 觏� f�<IR80� �|42� ef��  @ ���~�N��� �� �|� �^ .���`��(��Z� �<=uD������ �u6;�r2�?��|�-u��� r�u;�r
�������ef��   ��ef��   fa�fSfPf3�f3۬
�t4��
�ufX��f������+<0r<9w,0f�f��   �u
gf��f���fX��f�����f[�SQ3��
�t13�3ҹ ��
�t$<Ar
<Fw,A
�
<0r<9w,0���Ã� �����Y[�W�>8��_�e�>	� .�>A u.�A ��e�	 e�	e�	 .�>�t2e�	.�>=t.�?  .�>>t.�A �e� Qe�  : ��X�: e�� e�
 $�f3�.f�G.f�C.�K.�M.f�>��tF�-�
f��
.f��f+��� .f�Af;�s"=@ �� %��ef�� .�A.;?� .�?f3�.f�?�tf��
� f��� �;,r.f�Cf��
.�M� f% ���f�u.f�?f��
f�   f% ���f�tr��+r�.f�Cf��
.�M.+?��f��
f�tVf% ���f�t*f�   ��+r�.f�Gf��
.�K.M=@ r!.;?s!.�M.K.�?.�Aef�� �ef��.�Ae��.�?e��� �.�У�� .�A���e��e��.�?���e��.�Уe��e�� ��e��.f�>У�� f��f> .f�6Cf��
f6$.f�M���3r!f�.f�6Gf��
f6$.f�K��3r�ef����fPfRe�
Af�-   ��f�г�X��f�fx+  f d  f�  f   fx  f��fZfX��>Z�uf�EISA.�>�&f;uef��ô���� &�G��
 ef��   �ef�>�   tef��   ue��@ �PSQVW���ef��   ua�@ �����% <uQ����d9 uE.�Ud� ��d� @ .�U3�3�� �f����� R�!���t&�_�3���\r
C�<Zu�D@��_^Y[X�WVQ.�>���� ���
 ef��   Y^_�P�$�p� � �q<1� <3�
 ef��   X�QRSP��W�e��
���!�� ����@ �( ���� =���0 ��f�E
ef��df�*�O�  f���0f�E�׹ � =���m � �*�q ���tD�  f���0.f�5�
 �3� =��t%�0.;5u.f�>9 t.f�9ef��df�*��  f���0&f�L ef��df�*�. _��X[ZYø=�!� �ظ D�!� �@u� >�!���Ã��t� >�!øD�!� ;�t���øD�!� ;�t����P��� ��  �؁& �.�>W��
 .�>Y�� ��.�&[.�W&�&�G��&�G�3����� t	f��&f�@ � 	tdf�3f�t&f�D �X��� �    SP.��*&�?EI�k &�SA�a � C�/<��V �C�/.��*.��*&�> Co� &�> mp� &�>  aq�& � .��*= � ��P�	 .�>�*t�.��*X[ô�� ��� ��$<� ���ô0�!.�`<
s<r	w��
r����.�>�t.�>�t	e�>	�uú��ʃ�����8� �t�.)U��3��� �؋��3���d�� d�.d�>B � ud�B d�>F � ud�F f3����� �ÿ�
�������&��.�>b�e�� �!�� �� � ���S&�>$�R�1 &�&%�r.�r �.�t���&�+�&�*����H.�r.�tQR����� ��p� �����8 ��p�1 &�&%�r.�h �.�j���&�.�&�-����H.�h.�jZY[�WVQ.�>���� ��Y^_� .���                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  �fpz(���&�                                                                                                                                                                                                                                                                                                                                f`�.��>u�t�(���&��3���� -�t���(�&���� %���>��!��ef��   t���ef��   � ��	�U �~ � �3۹	 .���>������M �6X�fRf��   �
fBf���   r�fZ���b�A��.�s��fa�P�>���cs�F=��v�X�P�>����s�0=��v�X�P� ��:s#�r.�>X.�X.ǅX �H.��Z���X�.�>��� �3�� �`�� `� r?� ��؎�3�� �� 0���� 3��޹� ��ح���= �r= �s��� t= ��s ��3��޹� ��ح���= �r
= �s�D� ����/�؋����= �r	= �s�� ��������= �r	= �s�� ���/.�>X.�X.ǅX �.ǅZ��a�3��޹� ���؋Э��Ё� �r�� �s��� t��&�?�u!&��u�Ѳ � r�� r	��� r���ô�r��= �r�����= �� ���The IBM Personal Computer Basic.�>��o ef��   u%�5�!��= �uW�� uR� ��  �I��uE&�=BMu>� ���3���.�6B�u,QW�7B� �_Yu�.�>X.�X.ǅX �.ǅZ�����	uHh ��>�_90uV�>�_/uO�>�_/uH�>�_0uA�>�_7w:�>�_1w�>�_1w	r*�>�_6r#.�����ef��   t.����.�� ��VW.�>��~ � 
�<�u�$
�<�tn$������ ��� � &�$4&�d��:�uK��R�ò�� ���� Zef��   � &�& �BB�$���2�2�&�����������ز� ����_^�PSVW��3�.�>�te�>	te�>	t��.�?.��\.��t	��.���_^[X�PSR���؊T����t���' ��� r�;�w�� ��Z[X�SR�� �� ;�v�Z[�S��.��-�.�-[�fQf�   .g��-  <tU.g��-  t.g��-  �8.g��-  t4.g��-   t.g��-   �.g��-  t.g��-  sef���fY�e�>	tKe�>	tCe�>��u;.�� u2� ����t$�>��� ��� �s� ����t
- ;�s���e����='  e�>	�� e�>	�x e�>���n .�� ufe���>��;�s	e�����M����� .��-�t
ef��   .��-C��؁� ��f�   g�M='  ���'���'�����=' �ef��   ��e�>	�(e�>	�.��? u\�> ���@ +���
f�6='� �����u-�� u
.�>�� �؁���$�����g�u?'  ����'�F �6='� �8 e�>��te����� 3�.���.��C��f3�3ҹ .�6�sJ.���3���e�>��t��v�"�� ul�� t.� - ����g�u?'  ����'��؁����BF⫉='� f�   g�u?'  Ng�u?'  +�= u������e��� �ef�� @  ��e������>� +�3�.��-�u>.��-ue�>	� e�>	�
 .�>�� .��-u
9>u�>.��.FCⷋ�.�.Ã>8tCf�6='�>����3�3��- ����u����g�u?'  ����'��؁����F �Ӊ6='�PQR�ӋӋ�3���� .
�-. �-C��؃��ZYX�PQR3ҹ 3����� ���ZYX�S��+���.��-C��;�r�[���3ہ?U�u6f3�f3Ɋof��f�uf�   f�Ѭ�fIu�
�uf���؃�������� �����h �f3�h �3������f�u(f3��ށ>B  �u����;@ vh  ��������Q��3Ҏ�� ����.��- uF�� �� ��� A��Q�� �� �������� �������������� [;�u� =��v��،��u� �����Y��  fVfWfS�Ȏ�f�6�Nf3�gf�E���gf�E��= �� f3�fP��� � f�   �� � ��fB��gf�u� gf�M�fVg;t'gf�^
gf�vf��f���f^� ��fXf@f��r�� gf�m� fPfQfVf��f�   f�  f3�f3���f�Ȇ�
�t�"���
�fBfOu��f3��f;�sBf��gf�f3Ɋ�2�g�/f��f�fJf��   rf��   f+�rfBf��f�>-g�f@��f^fYfX�I�f3��f�   f[f_f^��fVfWfS�ȎرQ� ��Y�� ���� ��f3��ؾ�>��� g�F"�� g�F"@�� gf�vsfQf�	   gf�Ff%��� gf�^f��f��
f�fKf��f��f=   sBf���   r9f=�   sf��   f���   vf��   f+�rfCfQf�>-f��g�f@��fYg��tf��fIu�fY���<�t<�t�fY���<����#�f�   f[f_f^�f3���U�� ���=�.g��-  �� .g��-   �� f`��׎�f���� ���f��ώǍ>�.f����3�� �f������� f3�f�D�f���fPfX�f���&f;�� f��f�^ f�� f��f�^ f�� f��f��f�^ f�� f��f�^ f�� f������f��rXfaf`f���   r8f���   w/�ώǍ>�.������3�� �f��>�.g�r����3�� ��f�t5fa.g��-  �� ]�Å�tfaf`f���   rf���   w.��-u�fa.g��-  ���V�6Z��t��;�w���;�r�������^�WVQ.�>���� ��Y^_�.�>� �) PR� ���&�>��'u����t.�| �.�~��ZX�.�>� �: e�>��t2e�>� �|)e��� 3�����u ���e����ef��   �     PSRW� ���&�> ��= ��� &�=DE�� &�}LL�� &�}XB�� &�}IO�� &�}S�� ��&���=  �8 =  �� =��� &�}��&����0tՋ؃��������� tċ����&���% � &�=��&�E&�=�����.�>0M.�2M�  .�0M�� �r� K.�>X.�X.ǅX �.��Z���_Z[X�               AMERICAN MEGATRENDS INC07/07/9104/25/9105/05/9106/01/92 PSQRVW� ����3��0N&�%��a�
 ��z� ���G�� �1 �:�uہ�GN� ��3۾GN�< � ���� �� �������_^ZY[X�             ��         ���                 �������������  �   ��    ��    �      ���    � ����        ����p@          �      �      ��    ��pp                      ��������    ��    ���������� �       �������� �       �����������������         ��         ���         ���  ���O��       ������������N��       ������������N��       ������������B`       ����g       �����������������       �����������������    9 �����������������  �  �  �  �  �  �  �  �      �      �      �      �              ���   9 �����������������  �  �  �  �  �  �  �  �      �      �      �      �              �                                @  /W/W/WSWAWAWAWtWfTfPf���@R�Is�&@R��*��f�JRfH��f\�fQfRfVfWfS��rf3�f��f���u��f3��@R u4f�6\f�\�WfSg�^tg�}ZR  sMf;�sf��f[gf�v���1f�6\f�\�#fSg�^tg�}bR  sf;�sf��f[gf�6��f��f[��f��gf�F�q	@Rf��f���f_f^fZfY��@R t�/�f���t�@R t�+�@R t�W���fQfV����f3�f�6\f�\�gfFgf�6��f^fY�fPfSfQ����th  &��f�   f��f��
f�   fYf[fX�fPfSfQVW�>�[&�=�� ��[� �u@� ��[�u7f�   &f�. f��&�, f+Ë6\�\�f9\ufDf)Drw�J_^fYf[fX���fPfSfQVW�>�[��[� ��uV����&�&��  �tG&f�� �>&;� w7f��&�� &+� &� r"= �w&+� f��f��   f��f�   �_^fYf[fX�f`� �� �C�/�BR�DR� �BR�FR�HR��BRf���]�	���BR�tx����BR�tl��f��f��f��f����  f�f��   rf��f��
f�f;JRvf�JRf+���@R�f�6\f�\��g�V�BR�tgf�6���fa���fa�P� C�/<�X� ����f���t� ��F�fPfSfRfWf�\  f�   �Af��   f��
�  ��&��f_fZf[fX�fPfSfRWf�\  f�   �f��  � f���>�[�ǿ���&�=&+� �&� &� �_fZf[fX�f`fT�  �����&��f��f3�f�\  gf�O��� gf�7gf;Vu
gf�6���p�gf�V��m fPfSfWf�\  �xf_r8gf+$vf�f3�gf$f�  f% ���f��
��fRf����BRfZ�t �fRf���
�BRfZ�tf����f\fa�f���f\fa�PRfQfVf�6\f�\��
g�V�BRgf�6��f�6\f�\��
g�V�BRgf�6��f^fYZX�fR.gf��NR  �W fZ�fR.gf��NR  � fZ�fRf=   ~f�   �/ �	f�   � fZ�fRf=   ~f�   �\ �	f�   �� fZ�gf�^gf^f��f+�vf#�gf;^rf����+gf�^fKf#�f��f�gf+^gf;^vf3���	f��gf^��f��gf�^fKf#�f��f�gf+^gf;^rf3���$f��gf^f;�s��f��gf�^fKf#�f��f���fQfRgf�^gf^f��fIf��f#�f+�f;�rgf;^s6gf�^�,gf�VgfVf+�f��f+�gf;^sf��gf+^f;�s�f�����fZfY�fQfRgf�^f��fJf�f��f#�f��f+�f;�rgf;Vv8gf�^�.gf;Vvgf�^� f��gf+Nf��gfNf;�sf��f;�wf�����fZfY�fQfWf3�f3�gf�O�8gf�?gf;Wt���(gf�_�gf�?gf;Wugf�GgfG��f+��f_fY��f_fY�fPfQfVfWf�\  gf�O�gf�7gf�f;�t7�f����f�\  gf�O�gf�7gf�f;�t� f�����f_f^fYfX��f_f^fYfX�fPfSfQfVfW�� gf�^gf�Ngf�Ff�\  �f�\  gf�K�fgf�gf�CgfCgf+Fw���Lgf+FtrCfSf��gf�Cgf�^gf^�M f[gf�Fgf+Cwrf���[ f���gf�C�f_f^fYf[fX��f_fYf[fX�fWf�\  �Z f�\  �~ f_�fVfW�4 gf�^gf�Ngf�Ff�\  �\ f_f^�fWf�\  � f�\  �C f_�fWf�\  gf�7� f_�fPfSg� tgf�gf�Fg�g�Cg�O�f[fX��f[fX�fPfSf��gf�Fgf�f;�tgf9Cv�gf�Cg�g�Fg�0g�sg�Gf[fX�.��[��� �.��[��� �fVfWQ��f����  f��f���[  f�  ��� � Yf_f^�f`���؎�f���" f���% A��6�[������rfa�fa�fPS� ��fPS� ����[f�����[���[���[[fX�VDISK(d   �� �03COMPAQ                      �      �                  \\  \\  \D{�$\\            4\\            D\$\            T\4\            d\D\            t\T\            �\d\            �\t\            �\�\            �\�\            �\�\            �\�\            �\�\            �\�\            ]�\            ]�\            $]]            4]]            D]$]            T]4]            d]D]            t]T]            �]d]            �]t]            �]�]            �]�]            �]�]            �]�]            �]�]            �]�]            ^�]            ^�]            $^^            4^^            D^$^            T^4^            d^D^            t^T^            �^d^            �^t^            �^�^            �^�^            �^�^            �^�^            �^�^            �^�^            _�^            _�^            $__            4__            D_$_            T_4_            d_D_            t_T_            �_d_            �_t_            �_�_            �_�_            �_�_            �_�_            �_�_            �_�_            `�_            `�_            $``            4``            D`$`            T`4`            d`D`            t`T`            �`d`            �`t`            �`�`            �`�`            �`�`            �`�`            �`�`            �`�`            a�`            a�`            $aa            4aa            Da$a            Ta4a            daDa            taTa            �ada            �ata            �a�a            �a�a            �a�a            �a�a            �a�a            �a�a            b�a            b�a            $bb            4bb            Db$b            Tb4b            dbDb            tbTb            �bdb            �btb            �b�b            �b�b            �b�b            �b�b            �b�b            �b�b            c�b            c�b            $cc            4cc            Dc$c            Tc4c            dcDc            tcTc            �cdc            �ctc            �c�c            �c�c            �c�c            �c�c            �c�c            �c�c            d�c            d�c            $dd            4dd            Dd$d            Td4d            ddDd            tdTd            �ddd            �dtd            �d�d            �d�d            �d�d            �d�d            �d�d            �d�d            e�d            e�d            $ee            4ee            De$e            Te4e            deDe            teTe            �ede            �ete            �e�e            �e�e            �e�e            �e�e            �e�e            �e�e            f�e            f�e            $ff            4ff            Df$f            Tf4f            dfDf            tfTf            �fdf            �ftf            �f�f            �f�f            �f�f            �f�f            �f�f            �f�f            g�f            g�f            $gg            4gg            Dg$g            Tg4g            dgDg            tgTg            �gdg            �gtg            �g�g            �g�g            �g�g            �g�g            �g�g            �g�g            h�g            h�g            $hh            4hh            Dh$h            Th4h            dhDh            thTh            �hdh            �hth            �h�h            �h�h            �h�h            �h�h            �h�h            �h�h            i�h            i�h            $ii            4ii            Di$i            Ti4i            diDi            tiTi            �idi            �iti            �i�i            �i�i            �i�i            �i�i            �i�i            �i�i            j�i            j�i            $jj            4jj            Dj$j            Tj4j            djDj            tjTj            �jdj            �jtj            �j�j            �j�j            �j�j            �j�j            �j�j            �j�j            k�j            k�j            $kk            4kk            Dk$k            Tk4k            dkDk            tkTk            �kdk            �ktk            �k�k            �k�k            �k�k            �k�k            �k�k            �k�k            l�k            l�k            $ll            4ll            Dl$l            Tl4l            dlDl            tlTl            �ldl            �ltl            �l�l            �l�l            �l�l            �l�l            �l�l            �l�l            m�l            m�l            $mm            4mm            Dm$m            Tm4m            dmDm            tmTm            �mdm            �mtm            �m�m            �m�m            �m�m            �m�m            �m�m            �m�m            n�m            n�m            $nn            4nn            Dn$n            Tn4n            dnDn            tnTn            �ndn            �ntn            �n�n            �n�n            �n�n            �n�n            �n�n            �n�n            o�n            o�n            $oo            4oo            Do$o            To4o            doDo            toTo            �odo            �oto            �o�o            �o�o            �o�o            �o�o            �o�o            �o�o            p�o            p�o            $pp            4pp            Dp$p            Tp4p            dpDp            tpTp            �pdp            �ptp            �p�p            �p�p            �p�p            �p�p            �p�p            �p�p            q�p            q�p            $qq            4qq            Dq$q            Tq4q            dqDq            tqTq            �qdq            �qtq            �q�q            �q�q            �q�q            �q�q            �q�q            �q�q            r�q            r�q            $rr            4rr            Dr$r            Tr4r            drDr            trTr            �rdr            �rtr            �r�r            �r�r            �r�r            �r�r            �r�r            �r�r            s�r            s�r            $ss            4ss            Ds$s            Ts4s            dsDs            tsTs            �sds            �sts            �s�s            �s�s            �s�s            �s�s            �s�s            �s�s            t�s            t�s            $tt            4tt            Dt$t            Tt4t            dtDt            ttTt            �tdt            �ttt            �t�t            �t�t            �t�t            �t�t            �t�t            �t�t            u�t            u�t            $uu            4uu            Du$u            Tu4u            duDu            tuTu            �udu            �utu            �u�u            �u�u            �u�u            �u�u            �u�u            �u�u            v�u            v�u            $vv            4vv            Dv$v            Tv4v            dvDv            tvTv            �vdv            �vtv            �v�v            �v�v            �v�v            �v�v            �v�v            �v�v            w�v            w�v            $ww            4ww            Dw$w            Tw4w            dwDw            twTw            �wdw            �wtw            �w�w            �w�w            �w�w            �w�w            �w�w            �w�w            x�w            x�w            $xx            4xx            Dx$x            Tx4x            dxDx            txTx            �xdx            �xtx            �x�x            �x�x            �x�x            �x�x            �x�x            �x�x            y�x            y�x            $yy            4yy            Dy$y            Ty4y            dyDy            tyTy            �ydy            �yty            �y�y            �y�y            �y�y            �y�y            �y�y            �y�y            z�y            z�y            $zz            4zz            Dz$z            Tz4z            dzDz            tzTz            �zdz            �ztz            �z�z            �z�z            �z�z            �z�z            �z�z            �z�z            {�z            {�z            ${{            4{{            D{${            \4{                                                                                        ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������fPfSfRfVf� d  f�    �� f���H f�d{  ���� .gf�^ef�D	�:f�-   ��f�г�X��f�fx+  f�    f�P   f����� .gf�^ef�H	��2f�i   .gf�^f���  ef�P	�0 f���( �f��  f�    f�X   f���>�c .gf�^ef�L	f�   f�    f�   f���r<.gf�^ef�X	f�x  f�    f�   f����.gf�^ef�T	e�>	t��f^fZf[fX�f`f�d{  f��.gf�Fp+  .gf�F.gf�~f��f�p+  f�f��� f3���f��f��Xf3�f�p+  .gf���{  gf�Af�   �.�f�fC��uپp+�f�$f�D����f��f+�f�>�(�Ѓ�>�<+�e��&� &�E  �>8te�>	t&�E��f3�����:I��f�f��f3���f��f��Ѓ  f�   �:�����f�f��f+�f�>�(�Ѓf3��:���f�f��f3���f��f��Ѓ  f�   �:����`�f�f��f+�f�>�(�Ѓf������:���f�f��f3���f��f��Ѓ  f�   �:�����f�f�d{  � �f����f� ef����ؾ �  ����f�f�&��&��� ��f�f�&��&��fa�fPfSf[fS���r#f��   r�.gf�F.gf�^� .gf��f[fX�ef�����fQfW���f��f��fIf����  v&g�f��&gO&gf�Gf��&g�G&g�_f��&g�_&g�f���� t-f��f����  v&g�f��&gO&g�_&g�f��&g�_f��f_fY�fQfVfW.gf�N.gf�~.gf�6���rf_f^fY�f_f^fY�Q3�f3�f�6$�Xf�   f�   ���rf��.gf�<��{  fBQ� ��Yr��Y�ef�����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      �f`���	���d �G�@0e��C	ef��f����X  �f%�  f f�����&�&- �f�B�t��
f�    �f�f�(sef��fa�ø������x��� ���)��� ��� ���e���  ���H ���e���  ���� �����  ���P ��	�� ���X ��� �� ��� ��  ��  ���� �u�  �u�  ���� �d�� �d�  ���(�S�� �S�  ���0�B���B�  ���� �13Ұ��  ����"&�G��f`���ظ���e�>	 u�>8t�>+<&�У�0�f��
&f�>��t&f��f+���f= �  w.;Av&f�A��&У��� ������
��
�Bf�,f����? f���� Ë�f��f�   �Ѫ��f� f��   �]�fS����J&�&�\f��&�\&�D�&�D�&�|f[f�   ���f�f�$�� ��O&�<&�\f��&�\&�D�&�D�&�|�����Ѓf�$g ���f�f   ��f3���f��f��Ѓ  f�> � �����Ѓf�<f��f��ge�>	���>8t &�У��'&�>. �f`.f�.f��.g8�.  t���� fP��~f�� @  f��   襪f;�fX�� f��f��f� @  f�   虩�� .gf��Σ  .gf��ң  .gf��֣  .gf��ڣ  .gf��ң     .gf��֣      .gf��ڣ   0  fWf��f� @  ���f_f��f��gf�%��f   f�f   f�f   f�fa��f @  I���-.gƁ.   ef��   fa��0u f�%��f   I���f3�� &+Уf���f3���f��f��Ѓ  f�> f�� 0  � �c��Kf3���f��f��Г  f�> f�� 0  �BI�Qf�   f��   �*��Y��f�g   f�$� �Ѓe�>	�� �>8�w f�6<f����gf;��c &�6У��X +�fPfQ&�>. t2.f�.f��.g8�.  t���.gf��Σ  g f�f��fYfX�fYgf�$f��fXf�f   Nu�f=g  u�us+�f   f�f   Nu�f-   f=g  �� &�>. �� f`.f�.f��.g8�.  t��� fP�|f��   e�>	tf��   �9�f;�fXr]f��f��f�   f�   �/�rEf��g fVf��.��-f^uf3���f��f��Г  �%��fWf��f�   軯f_f�fa���g.gƁ.   ef��   faf=   r$f=   s@f-   ef�f�f   ef+��&fVf��f��.��- t e��f�%��f^�f^f�f   I�L�f3���f��f��Ѓ  f��f��   � ��rJ����ef��fa�e�� t@fP��� ��e��3���f�@ ef��df�/��f���7f�@ ����e�6����fX��e� 	t3������ ��f���<f�D df�3��fPfS.�>�uE��zf�� �  f��   e�>	tf��   苦f;�r"f�   f�   芥ref��e�	f[fX�ef��   ���   S���&�&�W&�G&�g[�I���AÊ�������Q������Њ� Y�P�3�P��X� �u� pP��X� pt�����X�PS� ����&�>��3Cu7�&�>��Ft.&�>��Rt&&�>��Dt&�>��Bt� =  u�$� ��% = [X�P�� ��X˰�� #�t�B�$ #�t�. =B t����3��SP�: [#�t��d�[�SP�) [#�t��`�[�� #�t�`2�ø���Q����d����Y�Q����d����Yð� %P ��p� � �q��p� � ���q�PSQR�� 3�3Ҋ�����������.������/�����ZY[X�           PW������ �㫋«_X�P����ë�«X�&��؁��% �&�U�fSf��f������f[�fSf��f���������f[�          �&,28>DJPV\bhnt@FLRX^dj�ef��ef��f3��)��H f������� .g�u �  dgf���  dg���  �.g�u�  dgf��dg�D��F�ʍ df�d�����             fS.��.f��    ef��    f[�fSef�>�u�X&f�_ef��f[�f�d�l u/f�   葢f�hs
ef���� f��   r�f�f��   vb.f�Uf��f��fIf�f=   sf��   uf��   u� f��   uf��f����  f��  ��f+�f+�f�hf��.U�l�[ � �ef��   t3۹ 3�����t�t0eFF��ef��   t3۹ 3�����t0eF��( 3���~�t0eF����e�6�
��f3��
 Q�րʀ��r�ր���r��?
�t.:��� .����	df�6��F���ƈ�Y�.�����H��f�
   � g�M$  ��f�
   f�df��f��g�M$  ��= � ��dg��  f�df��f��g�M$  ����= � ��dg��  ���           $debugdd emm386     � @P� �  AP� � (@P	X   P AP))  AP)) AP��  P��  P�P   PeH    P��  P11  P`�Ȏغı� =�!� �ظ  �غ@�0�D�!�>�!�!�  �ظh5�!����� �C�h=��u~�@Yf�.�
�@.����B.�±��3���3��p�������G  �G �G��G��G �p�H� � D.��������ؿͱ�Ա� ��؁�  Q��ȭ�Э.���Y��a�            fPfS��� ��ef�H	f�)  df��f3�f�شR�!��f��f�f��"f��)f3���f��f  f��)�f[fX�PQVW��e�6�
�؎Ƌ��>B��� W�<� <
� < �	 < � ���&� _P�D� �� ��+�`�!X�D�_^YX�W����_�           `�3�3�.�.��.��.�t!.��-t�(�.��-u���Ӂ�� �FIu�e����� �ӎ�d C��d�  d Cd�>  u'<Zt�� ��d C� ��d�  d� d) d� ��<Zu����� R�!����� &�_���& r{C&�>  Zu�e;�uk��d� Cd�>  ZtC& ��& C���@ ��d� ef�� �  3�e����d Cd�>  Z��" �t��e��d Cd�>  t� ���a�fPf3�df�  df� df� df� fX�SQV�����3�.����t��:�u�;�s�ы�������t8;�vA�� u��.ǅ� ��.:��t��� �� .���;�u��� � �:�t	�Ӂ�� � ^Y[��t��d�  Md� d) d� �e����d�  Md�   d� d) d� d�  d�   df�     df�     ��d�  Zd� 
 d�   d�  d�   df� SM  df�     ���e��
r9�� �> �e� 	t2e��
s+�c+ ���t!�c+e�& 	�ef��    �
ef��   �SPQVW��� ��e��
e��
d�.�Y.�W&����� ����P &�w&�G����&����: &���1 ��3���.�[ �d�&��&�E8&�e��.�d.�>b�
ef��   �_^YX[�PS� h  &��
�г�ҳ��s
&f��   [Xôh  ��
ôh  ��
�t����S�
 ��[�S� [�Q�3�3�&����d�>  Mtd�>  Zu&d�>  ud d; sd� d Ad�>  Zu��Y�                            �������d��( ��� �S����S�� ��� �B����B��  ��� �1����1��  ���  � ����ؾ �������f�f�&�Ƿ&�ŷ� �ȷf�f�&�Ϸ&�ͷ�.�ط.�&ڷ�f.��f.ȷ �f��"��|� �  �؎��Ў��� �f%���"�ꚸ�.з.�ط.�&ڷ �"؝�              STSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTSTST                                                                                                                                                                                                                                                LE             �                       *   8      q       �                       *          5  M  k      l       �    *� 4                                                           E             ,                   *    @                             LoadHi    �        �  �  �       �D b�
 �� 0�
' 	` �F �
' LNx' 
 �� ^P �� Q� yT U ;�' # J �Q �X �X �� J� �� � [
' %� �\ Y� �  
' ��� R� �  +  �`' $6 �du�' $S �x �d' (? � �n �( �h �h' ��? Tl �� �0 h� �4 y� ��
 �8 � �; �< � �} �� �� �' @E ' a� �@ �   2� SC �
 _D i� �� � yE v A' H�� �� ^ 	' �b
� �
�' 	H��' 
Rkv~� 	� 1� �� N UO' 
� &�� � �� �P r� 1 �	�' ^}' 
���,2 ��' T`I	 �� �' 
����	 � �� �	X �	Y mY � H' *K' 9 X�' 
8 ' ���; �	\    �'  Z���$  � _	 ' `

 	 '  ^� �a' !�� /" _c' d9
?
hn �$ �� �� � h &	�' h]
� �(' (���:FW A) ��' ,@�' �	S� �� �� �� �	o ��' 0�� v� �' 4�� (�' �D
s Iu �x �x O8 ��' <�4 �| < �� � ='  � � ' � �' 05 O  � �' ��                                                                                                                                                                                                                                                                                                                                                                                                                      � �  VW�  �5
  Ftz3�j PPPPSj �5  � S  �� �t`�=$  �;�=(  �;���  ��
�5$  ��`   �	  ��   �< t�����RQj jj PjRS� `  ��YZfB���_^����� �  VW�=(  �4;�t@j V� X  ���u��`� 
  � �  a�� �  t��tj j PV� V  ���t���`�[
  � �  a��_^�� �  VW�   �=(  �4;�tUj V� X  ���u��`��
  � �  a�� �  t��th    j PV� W  ���u�`��
  � �  a����_^�� �  VW�  3��=(  �;�=$  �;�����tj P� U  ��_^�� �  �5
  F��   3�jVVVVVj�5  � S  �� ���   �$  �(  �   �QI���  ��	  �,Q�=$  :�r�J
�fJt���fJ���Y����YI���   w��   3�h�   PPPPSj �5  � S  �� �tL�5$  ��5(  ��5$  ���
  ������3�HÜ�`��
  � �  a�� �  t�����`�;  � �  a�� �  t��`3�� �  � �  �=
  G��   3ۜ`�}  � �  a��`��  � �  a��   �QI���  ��	  �oQ�r�J
�B���uF� �  ts�`��  � �  a��`��  � �  a��`��  � �  a��`��  � �  a�3ۜ`��  � �  a�CY���YI���   �p�����`��  � �  a��� �  �  �ȁ�   �?  �Ç��  ����P��PSQR�u�j VjR� a  ��ZY[X�����PSQRj jj VjQP� `  ��ZY[XPSQR����  j jQSR� ^  ��ZY[X �"ߋ}�Q���  ��	  �u��`��  � �  a�� �  t��tmf��@ QRQ�=$  �<8:�rs�J
�fJt���fJ���Y����ZYQ�5$  �432�z{�J
�fJt���fJ���Y����Y �"��Ü�`�   � �  a�� �  t��� /  Ü�`�U  � �  a�� �  t��� /  �� �  j�� �  j �<$ t4SP���   ;�X[u$��`��  � �  a�� �  t��`3�� �  �   ���   vI9��  u�SQ�   P������XY[���X�� �  `�H  arn�=<   te�� u�'  ��u��.  ��u�*�����u������u�J  ��u������u������u��   ��u�  ��u������� �  �  �   ��  �t3QPj jPSR� ^  ��XY�u��`�l  � �  a�� �  t��@���� �  SW�=T  �[P�t���  _[uS��+\$����   [s�%\  �~t��%X  � �  W�=`  �?�%d  � �  f�AY_�%h  � �  ������50  � �  �54  � �  �Ð��� �  f�}Xuf�}u�=L  �tf�M,f�E ����� �  ��lW�|$� �  _� �  �L  ����f�EX�P  f��� f�]�!   � �  �L      � �  V�t$� �  ^��l���    � �  ���  � �  ��=8   u3�3��þ�1  �   ��� �  �   �  ��9Es��%D  �   ��   � �  ��� �  ��+�  ���  ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          ����            _PageGetSizeAddr failed on INST handle _LoadHi_Resume_VM
 Couldn't lock Instance buffer _MMGR_Resume_VM
 _PageGetSizeAddr failed on INST handle _MMGR_Suspend_VM
 Couldn't unlock Instance buffer _MMGR_Suspend_VM
 Allocation failure LoadHi_Inst snap _LoadHi_InstanceInitComplete
 Allocation failure VM1 LoadHi_Inst _LoadHi_InstanceInitComplete
   Start     Length
  
  
  
   Start     Length
  
 #ESI   #EAX
 No Instance data in UMBs
 Non-Zero flags _AddLoadHi_InstanceItem
 _AddLoadHi_InstanceItem bad InstType #eax in #edx
 _AddLoadHi_InstanceItem Links not 0 #edx
 Missed head detection _AddLoadHi_InstanceItem
 _AddLoadHi_InstanceItem LoadHi_Instance above MAX_INST_PAGES not supported #edx
 _LoadHi_InstanceInitComplete no instance list
 _LoadHi_InstanceInitComplete entry is 0 size #esi
 _LoadHi_InstanceInitComplete entry is 0 size #edi
 _LoadHi_InstanceInitComplete entries not sorted #esi > #edi
 Odd Case, instance overlap #esi @#EAX len #ECX
                            #edi @#EAX len #ECX
 IIC new Page #ecx out of range
 IIC Starting new Page #ecx, table struct not empty
 IIC adjusted inst rec to 0 or neg size #esi
 IIC overflowing size count page #ecx
 Computed LoadHi_Inst_VM_Buf_Size of 0 _LoadHi_InstanceInitComplete
 _LoadHi_InstanceInitComplete Temp_VM_Data_Area outstanding
 Allocation failure VM1 LoadHi_Inst _LoadHi_InstanceInitComplete
 Allocation failure LoadHi_Inst snap _LoadHi_InstanceInitComplete
 Allocation failure LoadHi_Inst Descrip _LoadHi_InstanceInitComplete
 Fail grow LoadHi_Instance desc buff AllocateLoadHi_InstanceMapStruc
                                                                                                                                                                                                                                                                                                                                                                                                 LoadHi_Instance fault on page with 0 IMT_LoadHi_Inst_Map_Size
 ERROR:  LoadHi_Instance fault on non-instance page
 Got an instance page fault on #ecx >= MAX_INST_PAGES in a VM
 FATAL ERROR:  LoadHi_Instance_VMDestroy called with EBX = Cur_VM_Handle
   �           LoadHi      �                      �                                     ����                                            LoadHi:PhysIntoV86 fails to map phys page number #EDX into page number #EAX
 Couldn't patch V86MMGR 1
 Couldn't patch V86MMGR 1a
 Did not find patch instruction 1 LH_Sys_Critical_Init
 Did not find patch instruction 2 LH_Sys_Critical_Init
 Couldn't patch V86MMGR 2
 Couldn't patch V86MMGR 2a
 Did not find patch instruction 3 LH_Sys_Critical_Init
 Did not find patch instruction 4 LH_Sys_Critical_Init
 Did not find patch instruction 5 LH_Sys_Critical_Init
 Did not find patch instruction 6 LH_Sys_Critical_Init
 Did not find patch instruction 7 LH_Sys_Critical_Init
 Did not find patch instruction 8 LH_Sys_Critical_Init
 Did not find patch instruction 9 LH_Sys_Critical_Init
 Did not find patch instruction 10 LH_Sys_Critical_Init
 Did not find patch instruction 11 LH_Sys_Critical_Init
 Did not find patch instruction 12 LH_Sys_Critical_Init
 Did not find patch instruction 9 LH_Sys_Critical_Init
 Did not find patch instruction 10 LH_Sys_Critical_Init
 Did not find patch instruction 11 LH_Sys_Critical_Init
 Did not find patch instruction 12 LH_Sys_Critical_Init
 Did not find patch instruction 13 LH_Sys_Critical_Init
 Did not find patch instruction 14 LH_Sys_Critical_Init
 Did not find patch instruction 15 LH_Sys_Critical_Init
 LoadHi: First UMB page is #EAX, this is unacceptable
 LoadHi: Allocate_Device_CB_Area fails to allocate 8 bytes
 LoadHi: Hook_Device_Service fails to hook AddInstanceItem
 LoadHi: Hook_Device_Service fails to hook TestGlobalV86Mem
 LoadHi: Hook_Device_Service fails to hook DOSMGR_Instance_Device
 LoadHi: Assign_Device_V86_Pages fails on page number #EAX
 LoadHi: Hook_V86_Page fails on page number #EAX
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           � �  �   VWS�} t��`��  � �  a�� �  t���U�B��;  s
[_^��%@  �B=   t)=   t"��`�	  � �  a�� �  t���B   3�9u9Bt��`�=  � �  a�� �  t���B=   ��   =  
 ��   B=   ��   ������5
  ;�tL�B;FvD�;�t5��;Fw�2�ʇN���u��`�h  � �  a�� �  t����J��r����
  �Z�2FtN�V�=
   t0�,  3��`   �`   ��	  �   j P� U  ���+   3�H�[_^�������`��  � �  a�� �  t��3���� �  �  �E�   �5
  Fu�`��  � �  a��U  N�>G��   O�F;Gus�F��^�O��W;�w��`�  � �  a�� �  t��;�w��`�N  � �  a�� �  t��;�v��`��  � �  a�� �  t��;�tSw���t���PQ�F�N�`��  � �  a��G�O�`��  � �  a�YX;�t;�s+ЉV��G;Fv�F��GF����t�p�����3�j	PPPPPjj� S  �� ���  �
     
  �
  �  �   �5
  �~��FN�N�M��N�M�M���]�K����;�tM��   r��`�"  � �  a�� �  t����	   t��`�C  � �  a�� �  t���M���;ˋM��]�t2����C���]�+�)]�w��`�x  � �  a�� �  t���M���  �B �J����	  �u��`��  � �  a�� �  t����	  �u�s���  ��ry�BtR�B�����؋�+ȃ�r_�B
+�f�Z�
  �ك�����;�tw	˃�+��+�ˉ
�B��B
�3���
  ������
f�Z�3ۈZ
�
  ��Z
�
  �

  3�f�Z�u� �}����6F�g����
  �  ���u��`��  � �  a�� �  t���  �=  �,  ��	  �`   3�8t>��B���   ��3۹   ��  �I��	   u���u����   w��
  ����3�H�Ü�`�  � �  a�� �  t��`3�� �  ��`�O  � �  a�� �  t���8��`��  � �  a�� �  t�����`��  � �  a�� �  t��`3�� �  � �  VWSQ�
  ��;
  v`�  )
  )
  j �5   � X  ���tT@jP�5   � T  ���t=�
     
  
  �  �   돋
  �
  ��+  Y[_^Ü�`�  � �  a�� �  t��`3�� �  � �  `3��    =
  r
�<      =   ��  �  ������ �  s��`��  � �  a�� �  t���`  V�  � �  ^s��`��  � �  a�� �  t���0  ��  �<f�u�|tO��  �<f�t��`��  � �  a�� �  t��u7�|t��`�)  � �  a�� �  t��u�T�c0  +���L�  ������ �  s��`�a  � �  a�� �  t����  V�  � �  ^s��`�|  � �  a�� �  t���V  ��'  �<8Cuu�|HtO�$?  �<8Cut��`��  � �  a�� �  t��u+�|Ht��`��  � �  a�� �  t��uf�D����  f�<�5��   �|�E��   �T�T  ��&  �<��~t��`�  � �  a�� �  t����  f�|t��`�@  � �  a�� �  t���t  �|tt��`�x  � �  a�� �  t���L  ��   �t)  f�<�5t��`��  � �  a�� �  t����   �|�Et��`��  � �  a�� �  t����   �T�T  ��=  �<��~t��`�   � �  a�� �  t��uzf�|t��`�Y  � �  a�� �  t��uT�|tt��`��  � �  a�� �  t��u0�T�X  �Lʉ\  �T�o  +��D�L�D���  f�<�=��   �|�
Q��   �L�`  �|.��f��   �|2�AYux�T�d  �d  ��  +���L�D��T6�h  ��  +��D1�L2��  �<��A�&  �|�  �|�B�  �D�DF�  ��#  f�<�=t��`��  � �  a�� �  t����   �|�
Qt��`�  � �  a�� �  t����   �L�`  ���   ��ft��`�<  � �  a�� �  t��uq���   �AYt��`�u  � �  a�� �  t��uG�T�d  �d  ��  +���L�D����   �h  ��  +�Ƅ�   鉌�   �$  �<��At��`��  � �  a�� �  t��u]�|�Bt��`��  � �  a�� �  t��u6�|'�Bt��`�   � �  a�� �  t��u�D�DF�D)Fa�=<   ��  j h�  R� l  �����!  �  �   =�   s ��`�Y  � �  a�� �  t���  �   �   � �  �50  �   �   � �  �54  j j� �  ���u ��`��  � �  a�� �  t���@  �$  ���(  ��  �    � �  s ��`��  � �  a�� �  t���  �5@  �_  ��  � �  s ��`�  � �  a�� �  t����   �5D  �  ��/  � �  s ��`�E  � �  a�� �  t���   �5H  �  �   �M����tg�   QPj j jP� r  ���XuY��`��  � �  a�� �  t���=P��  � q  XYs��`��  � �  a�� �  t���@��   ������`��1  3�� �  � �  =�   r=�   w�� t
�8  ������ �  ��lW�|$� �  _� �  f�EX�!   � �  �E�P  f�EXf�E  �!   � �  � �  V�t$� �  ^��l�!   �  � A  �!2  3�3�� �  �(2  rI�3��(2  �!2  � �  �(2  r,�50  � �  � �  ����   ��
�t���뿰 �빿2  3�3�� �  �(2  rV�3��(2  �2  � �  �(2  r9�2  �    ��G��   ��
�t����2  �   r��  r��Q   ��  �? t"���  ����%��  ��G�(   ������� �  �Y   r��   r�   ���%H  � �  `���54  � �  � �  �     �@    �P�x�@   j P� �  ��a�� �  VWQ���50  � �  t����   �t�50  � �  u����Y_^�� �  f��uf��  � �  ��   ����  �����  ����  �   +��� �  WQS�=   �������߃��3�f�G �tVW�
�   ��_^t$�ڋ?��f�����   �ρ���  ��������á�  ��;���   ���?Du5�GH��;�u)SR����;�Z[t�G���W�l;�wk���׋�+��]SR����;�Z[t�����R��;�Zu�?�ρ���  ��������܃��?Du#�GH��;�u�G����+���������[Y_�� �  �=  �  (C) Copyright MICROSOFT Corp., 1990 LoadHi  LoadHi:Sys_Critical_Init Fails         LOCAL GLOBAL                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         �� u�� u	3�3����=
s� ø �3�3��  �#Win386 LoadHi Device  (Version 1.0)  
LoadHi_DDB                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    MZ� :   ���*    ��R   !PKLITE Copr. 1990-92 PKWARE Inc. All Rights Reserved   �p      ��2�    �                  ���"  ; r�	��!� Not enough memory$-  ��-% ���P�#3�W�D��ː���S��9 ڌ͋���������Ƌ���NN��+�+؎Ŏ�� ����u����� 3���� �8�����A����B����H����M����S����g����h����i���r���Jt�s�3�3���Jt�����Jt��Ӏ�s(��Jt��Ӆ�t��Jt��Ӏ�r��Jt��Ӏ�w}.��	��3ۃ�t*��Jt�r#��Jt�����Jt�����Ju����Ӏ�s.��/���V��+��^�u���Ju����Ӏ�r���Ju����Ӏ�r���Ju����Ӂ�� ��뻀���Ju����Ӏ�r��Ju����Ӏ�wE.����t�Z��Ȁ� <�s�M�P�� �����  ����Î��؋ރ���Î�X<�t)�������Ju����Ӏ�r��Ju�����.�����[���3�����Î���&����Ò���ҋ����S�P�Ŏ�3��؋ȋЋ�����      	
                    	
      z U��  ��tV� P��M  ����G��\h
�u���>��
4�v���Ni% c!�>*[ t
� D/
�
�
�D
�
�X
/e�
X(� �^��]#A�����U�O~+�P1��U]�F����^�Ƈj]��~�r��\5t�m#D<o �S�u�E�F���a�Ae�
et�.�U�] a	� 7�sms�U�g���u�uKI��u!A��u������ ��g��*ſ���[  ��Q��@��*�;��'w�U��  �oX�`���/00k �/:�Uu'��;��u l�f�f�w+x������<�����+��v�X\���l��)� "��<�D�us��=Q#㕍e�/�SW$!z<IM�G�  F���n����9�R���w��L���P�6���Qkt�F��4��E�2v�|@��T�y���ɐ��}*��PK�h��R9��t�RX��JJw�F��:�����j�5�r��h��\RQ0	�m<�nK�uX>�X�u�fXQ�V��^���r]Y/��O\��!�ɔ*�=�*�#6�2�J���&�!!�Ap�3^��]Ð v�
 �qVƉb%h)~j�]3��'�L�x~^���t��p����98r���E�z����R���R�,�U�L-Lu �~���:�1�R�1�)TT舣-��gɈƉf�0�.#�&6�X�X]Λ+
��Oܛ��Ah���]�7y�+��۸. �f���1�(�������y��7t	#ܜ~pr����Oxo�:oM�Q���Q�+Q�vy��Ň�������Zh]	8�ڬ0 A�F��=ai$�=1c=2�a=3m=4=5  �2+���s�������' ����G�<@���f� a�S�Sb��H}� �� �o��H�UP���3 3+�T,�*��4+��)݀)�AΎ����Cg����*����7���
7�**v7yh�AW��W/U8UUf<�U� X$� ��)���6]�rL�MGdL�GVt�� ���Bm��O$E���S� �n"4sz'j�4�N��4�4�S�l��3�K3�yM���[ʝ9�9. R%,T�3��K+�Ug	�0+x��+6+4+=
�n�S�.)Ji�1�5
K-��/ ��l/�n�/&{�RHH�(o�/�("���'P8�O�6�������Z�BߘZ9V��$�2�2�(%�
q  ��*�4"|�.|��y�*
u��~�k�s2( ��F� ,٨<t<t0<u����8�B%�"���>͕
��\�8z���#���'�B��HH��,�<P�`�-0 l��� ��(�^�.��)�$����Θ�k�&�89��u�(��&�t�H�����ԧ� �F���6�4D��<��P���3D^�~즺 PSS�fȁ�����Q��}>�us��92P0P�&�����Z���-����)tk=�N qta�\�v�Z�"�QE6PFR�G1��!��[v`t`�`�`��.�!&�o�$T��}
0�
�

�躐&��K6� �'j}�W�`8o&A"l �l &���
&��%H��5*H�H��}���$�+�I9���&g$g���%3�,3�3��  6
6w�D%�N�r�~ ,r��y��������5�v�V�uP�!p�4V��{J�z71~x~;~� dV�~�r������t��-�H&:A^_ Mb ��h�tM���Ql*mN(N�$1;��k8�  ���H�N�*����N���vZ~�r�~�	6���F�%�� ��$�v��`����D�oD��������}(�8Q��#����&��C>��h�N 	�L|�����6$9�2 �q����� �W7sNK�����|��t��(��+u)�	�|���D����H1E����.,S��#	dm&x���H�e)���G4T�P=�t��A.�q/b����!��u�
����F�4�P;��!n��(8��]u"�*>���>�����?�Rj�� ̀���I'�2HFLIJ�"T�J���Js/J��L]RRDP���ț/Q���K��]Q�yKG���F�t@&��0����a����S�: �C�G�2T�cXR�Ȝz�ȓ	�	� ��LZ�\+�A�V������"�L�)��D�&}�����,�g� �!� m�v����B���i\����- �-�L�V�v-��ё�|S�l~S��V�� �-���
 ��0�^���&���n���T�#�# mC�S[�;!,D�B/B�Q�z�u�3^|�]��$���'���Z��!8@����)����y�s�w#�w� �(�)Kc�i��	��00��5�=�5p�����C�~,�>8�n���8�H�
��V�L*Ӧ¦|Ȅ^�� 4��apE��C���S��$�QERR���u((]�.E� ��c����I:h8����X�f"��D2/}W_T(mĈwNG_r�b�?�+��u��otp�<�4����HK�%$��� U����2DK�Q�����������S���2p���.�{�E�w<t`�� ބ�u%FT`W�@`M�H�v�	`kI�M�-Ј�qC�D`�`�`,`p8�&�����8`��nA C[�L����a�8J$?Т��R�����Am �ܫ������N��21����%��q�U%��ň(�^"�B�<3u<��?T8�7����*�(T�-�-��.JB>�|%�0�y�#?�5^�FhCtiB@
@
�@��Z�j �UH[�7?��;)?)�;���9�~��S�{�y���	� �%boP\�A|� �_`V�7���A����R��U�As?�1L���C�����oN���^N��H\Z�4;��x����  ���X��4�*�+�QP����L��wR7�  w�F��V��ur=@ �Ds���!$����]�
� ���J�r�6��=�e�=e�,���@����lnm? �4&B8r�R�̠�~�~ !)H@�#M
%ȚT�c�
9@�;�R��
��M�R��8Ҥ���!��Ѡ� �p����ZMr3�6M_+�A��>;A�$���Wu��K�!^ɵ�?� �O�S�Q�=ZZO�W�@�W����);Ƈ�?�S���x"6���]V�c7w�Fx?x�F�x�(�x����G))��Z�q6�#m+�O2$�؃�RI7��W�)`E_*EIEl���T���=�f+4q�4��+�+�c+؋�'��A��v��s)�2]�F+2�2�]6�=�S��� pstA�|�mNUz�*��=B@�jt��~��vF�tep*]O���Mu�>2�(+�3oW���*st�#�U�,aǣג�#d�T�p,Vx'R������<���'|�J;��l!>�-D=��� �7 �Da�J �Y�[IY�<O�ܬH� o�Yn�RY`[2��&�-(�-�9JT-�)Q-%$��JE-x9I����/�#��L!w�
Ttu����y��+�n����PI�+�n����+d������^��l��~4uQ�� ��)�bJ��Fb�b4��� ��� R�� ;���:��H��T��MR�r�d���;Ȼ�:��$��S�I>"�*��, �%����	K
�SH���/s� ���X�-�i�V<�R��F���tH�(�F�9�������Wq���ڜ�6��66���6���*����8 &q���%����U��Іwf�8<
\E01��/�7>kɔ���U���Ą|�+�w�@./�/6����&z��͐;�6
Ҁ�~�k6��@�"v�`DI
�*�koL�*�T*���1����Mt	�B	��r	�aA����a� ���6���L��A��� j�8�2�:�95����I$v��Q�!�j�&Bt/OA�W �s�g�n^;q.x!�Mj<�$�]7����zS����S�E�Su�$��-0�7"%�%�j��J%�#(7K"C���()���3"d���D�m6f ���uU�s��%R� }��R�os�Y������ �H�Z/� �z������#t��u�{������&^���V4׽�r�fE1��/{�͉�����<Pډֻ���Bː�ue@.�UsUS. �ݞ֗2�ϞtȚoޞܞe�`��-�5-��\�:@u� T�(m�N&��Q����r�o$���M�t�X1YMh�C?�H���q�,0�M?I/�4�d("��� �D�񃖁��k	s���������Rx�� ���B;Ư/��}�BC}Ӻ-1 �����;�u��#v��t�t������v�v�Mo
Ƅ�� e�C��Et0$y"�.�2Lh��]�3��2ׂ׀S�&�T~f8������J�@��T�c���5�$ �Q��R#�8h:BH@S��&L"#6��Y/ܤ�Abb	-d>�X0s^��1K��%�1FtD�t�Qk��V�v ��f�T�|�����2堿hQwR�2�o�JuHucu&F!o�� 0Uv�� ]ve m��(�;��r3��l��P��Zo�<�i�/O�d@�>Ht'��Z@t >�e����&j�6ƘD�.T��"w5�P@0I[C;n�*6�c�gE���L"��W*�=(	O�y:�Uu,;pz��u%�} ��<��v���� ���	�戀���ۑ�r�n%���O�X��H(v���� ����f�������t�y�u�$�?
v
8%� ���������{�w�+y諒z��V3{
3���1|À�+ұ�g~����������K���'��Ԋ�*�&���KgK�K�W��KV�#��ep��� h�~����f�3�E�ļ$f���0���R���U6�7)�U�)��)�)؊�����oKKƄp$�� �>tS@~�~� ub�k�&�z�5�9��"R�Ǟ�L
ƀ���~���t���?�t)���f��l�I[;��w�x�u��!a'��V�@L�=S���3�bOw�bW���u���5\����W�	�>�yn����S���
ʜ]�����saA�*:�t��ʙJ+��Xm��6e��ƅtgѰuvǅw��|z�{|`�߅�]��{����]DK%�*��&��F6�]��_4��v�S.�9��n!8�dJ\��%,c��� �� C�w��.��X��\<	܃��"9��dC����@�U��g�z[0 m�!�Ճ	�ّ�t��u�
�+�#��u� d �J;,o}��k7ku!\?k�k Ir9���%��2�-H�RKVPz��zC*���/�)�w^�ƀ��/�_���9%�jN%	%��M,p�F��D�!�v(��B��}N��sM�G�]�;w�&�RLF���AV�q=���X t!�@%���r�S�Pʏ=�lã��Q�^c�k'\����� $�����v�� PG��ۃP�;��ѧ��� O�'DO�\�-� mw�"� � �IWV���d���
Z&�{ɚ $)�B줄�*�%�$�p0+�+]��F�P�z\H�+�w� ��SS��/]/E&/E_�@/�</�J�~�h/�/��A�t���+k�w��a� �7]7]27� 77]P�C���S�� A	WZ[�S;� y8��"��Z.�s�	D_��,@��ZD��Y���3t"���T �ZO/*g*�WV<2Y� �g���w]�� ��F�~��������� t��t}�!� �����t]�^���\u����"�v��%�C$,X�w��Y'y^N�z �Tm?{%�?�=|)"�gK;#_Δ�����J���m.�ʳ	�W�^Wsr����W�W��2+.jO�&��] d]@P�0@Q�{]d�>�%���&M"K��p����v+�0�Q�)NpN�]X ��*3v�~�>��0_��7caCPVJH�v�P~�B1o��駁��32s] A��r�)��)	)mo|%�y�AxG�I���]�-EV*�8k&H�r]� �/�ZR�ĸ�PLU	"���p��ZC ���^�&�@ BRAtX�F�����0��]}$���KbB�Ȝo�8��u܊L���-�*�s����;�\�UrJ��p�n��
lS�`v��X�d&@����t&��"�"��"�"EN"�tQ�}a^��^�u�&DׁS@T�7 ,�P�] a  	ø@ ���r 4�5�t�!���t  } �SO��  ���}R� C���nV��$� �)�^&�?�^o�>q<�q����܁�>D�rB�����2��T��"��=��`=< tH1�./$���/���v�b������q"v���� i	)� �c��3siIaFrn~;�!�-rB?=C�@H�-I�u�$�)�H
#������߀N���&6f 6����P�x��� hݠ� "���q�F���	�L	.��:��%
'�ZP/gw��h�]���Z�Y��>+9!},#?�D ��7�/=N t�=O �4
�=R0D��=S�=W��YA�j�16��X�<>l`�������Z��qVt!�^ ��
&�/-���V�!!u]2�Eč�(-0 �'t ��v �O�G�3.����]��
39X�\��z�1�@�P�?�4�QQ?4�|�=  d`���P�F�P��Tװ1����(��
�
S&7
�
T
�
Z�U�Cn�:C C�o"C&+@;0��v ���ƀ; �����r��`�s�R�RDV^JZ��^8Vi�W�iX�MY��W��?�g�X�4MZ	[�4
\a���>VPōF��F�V��s���~ t8 �vA�
��^	^�F�2��$t�&� _�"ń�Nw9��2CBP��9ҍB=	3bII<��������� J�0 ;�s}�K�O�0� ���c���00��*nt�
��� Z��at��^|,�0t�@#�� ,�pta�S�1T�-9q�T�U��sH��S�<�%!�%|:T��^a�x�O*NFNu�� u��r���6b|�����<�6��ZВ���h�G7���Z �7�7���_�7%Rg�%���7	l�L�x۩���������$��bOD���lZ �q-��@�ZN���N�K!����o���	o�Z�o#q;�����n��ֻ�R�mT؋�Viq�>���P5� 5QQ ;dm�����=��~z��Hn{1�*c=Cty�x�!$=�����	�9���^��p��F��1�9w�8 0HW�v��`�#��.�99��>9u�����j�[���
����+���3��kP6�B'YN�;�5�� k3�T�v=�U�=V�9��9 9?�Q�
�dK��,��aJf�^?e=SN��s6l0�Il 0�ȉNZQ�7���"-L���1E���"� T�Ǣ�r�㣉
�%0@�=S|=9 r�v�r�r� �0U�9!߀��"�,9V���]�sC��u&�b4� T
#Gu\��V�@8#":Fm� ��-��3��`w�
#w�w� ʅ�3hL��t�q8|�4�lZYz�ɮt!UAa�S��L,$���-Ah�@v��IyL��ie��Ue�B3~7�d��Z�zL�ѓ.|u�TR��&eG7@��V��䅋V
�D��V��7^P�<��P�*��7����[쫤_s�*!��^�W�Ŧ½�KjC<��u#} ;�ɞ]T�b� 
?.J"xUJg��1SJl&�
��'����(��w,��N�ُN��p���0v ��V�F�V���+p�&�Gq��G���	�+�x� u˩ �wX�@PI�5�\��J �*�=G�=K0WV=Md�@t*� TQ���� ��� ԣ��@5� 5���5��5�����x0�1�����q�hM vv]�tau��	�z�cd��GE�&Q
Q�C�y����p���W��@jHuI@G;��2����G4V��S�j �%�+�=�����=.$G��p���q�ME�FT��MM�wH����< uW�T:唷��)P���S�GӾ��=������N�d
�
v�;��Q�APO�J`|뿡LT���H��N�P�Ra��T�@V�= t�=d4u�=��=�����V&���#�1 %���.���=�P�w_*W���}{�	��R�#��&���P;!/�6��1��{R���&��=)�!����P����a
��&$	�ؼR�3�q���S�����a�j6�
 T��Q2X��!� $_X�Xᢖ���*������S�I��(瑄�<�ӵ�N���O1��<r�?�lE�Z<�s�<�s/����&RH���qNm_l�q�	�� }[sM}�!�]����{��D-�]�3���J���]�:�sQ;��;[v2�ɵǺ��\4��u@qc�._�`u�Z``+`��Q�\�;�& 0WV��IID�����EC��I�:�E��$��'ё,d&��AQa�%�r�Zb�D�b��9i[^�h�'��؊��p�� 	hk�~�sgjO)�)����-�#�-��a]x�ha
�.
] �8XX���U��w�%��x
t�g��t~�.:]R���z�R��ȹp �����{�o�����r�\��M���	/b�)�t��#��T'і��S�1�F���� �j.��WV��]���6ЛA��p�/D8�+��u��KYN`L6oej
h�#j2�
 $��ܡ �������ﹸ����{s��B�U��d-(d���������Z�P�D%�y�$!�A�K������qC��N(N'�演�r6�66��,�~�s^�?6��D�<5u���)��c� �C��� 
+5�]������sH^3f�����s��`Ӿ�!��]�u�����B*�9�.D=H�`�Z��s���x/����  �n����Z;�`E��v��+��?�Z�� �R�PS��J��{o�VTJ�0B�7�ZX���{�^\���y�b#�`��'<�o)�� �@P�Pd$����?�7�f5d5qN�5
� >(�R�0���F��Ѕ�ۍx�H��X��$��ߥA���9S�ę8����,1��"Ըb&)r'
�X�+WV�$�	 � ��n���fR�L@ N��PRT�L|�#�"��\�|�J����+U"�d��[���u�V2�2 ��w��t�D����ޒ�+/���)Ջ��$>�R�/�YT���?<[Z��0�\
�$a�لx����vh���ڴ�����߀���4ɽn����|���p9ft332�+H��E��ڏ�%����t��3�4�(=�u�Ko2\$��_@���ۉOiO�W���#���R�^AQ	�+!y!T�J����L��3Y�_8����؋���t�%�����~�ٶ��d����N�E�
�=�V��jI�"F�NJ��"��`�P�9��H:	@��VP�"P��R�6	�߷�9v�s�P	�����+��'���pt>ʈ\h�˯�!qx���*�)���@�}!��_���,!��]!�n�Q�,��uk� >��yv\��`�
�5 U?�La���6��� �F�b!-��r
!Y�&�+3��s�5���2���|��]��"}⋼GB�#8P�#�ƋR�$��^�[�� 9r�����Ҝu�t�tvCI�AeǇ��F'�F�橾�:O�����|ҸO�<|k��6�:�U�䊔�:&������+� ҈�Ew�N/]������@��V�@�̵�j���%���τݓa�T�����ͺ�t픛D��ǉ؀��K�9���	��|]�H�^���H�A�=��2��	Z��H�*b!!���y����������(���e�=B˖��^���~(�+M�ǯ�
��=횥�t��Ӿ��ҩ:��U�ُ���9틅}+�,���j��m?����(��  �`*�����*���F��+'�6
�8P$*���?� ���n��J����+��E5U��hݥo�e�8J�����P� �V�؂� VA �Y"���t^7���i�NEy��#� ��w]��h9�s��u�y'��ł�!V'jp"{}"��&���X�ԩҀ�۰��D�S���W�C}� C�+��u�2�@B^�@25�@�:0�
�t�iW]�4��<�<t�>=R�� ��R!KR]������Y��]OB�B��s5I�UKހp���tGT.B}{�B ��ޟt@���@���@t��<��>0�w���7Z����x�e��.�|��k{LdҤL�)}3SvZ�8Pu��?������^jV^�o��)C�gh'hY
�\��կ\�$\���9���� u�r���]�v�z7\�GSP�Vس�Hn��v�Kv+�P�~��1�` ��X��J[� ��JÆ�t�(u
��GG bG�G[�#�
��ǩ�I�`-LT��\&ق%ߞVʛ5_�t�IխLRe���X8E�##���#�Ym�g��[WV���F�<�P��~�uInK���.Q�����;
Ƅ��� �	�yr��6���Lƀ,��� �y���0g��;^��r�F~ƅvy��4���{���X��z���n��6 u��{X`Q{�u���dF�"��Q*��wR�d�+���8�S4�����0E,+�Q4)�V������|H���^�ߚY=���?~�?�@�3iz@~@p����~
�����e�\�B�*���l@���+��5�0/��C+H��6�vD�'�	�w�/� *��yo�V�W��pc@B߳.�� �RY.0CS�{�P��
�9ȁ���Q�-�o%��!/>�!w!��� � 莄��j�5�嵹�T�)C7�t] 7�R]��R]*TR]R]�� j��X��!u!�]z��]3�c@+�r�02z�+�]qw];��~]ǅ��l�rw	
( �+r��d�]PC�]�6�3<󶲇�]�? ��]\�����Q���A<���� �ȉN��
+�j�� Fy�T�T�H��H ���]Q���+��ۓ!�!�+�Fڰ�
z�����V.*z��P�5uvǄ��yE�z{|;+������IO����t�	����MPK�L�����l�l /}�*!^�+u�23������]�v](��]��Hz{|]�ߖ]�����3�]�]M��%Phͅ�*��z=�P*>_����V�H���]�=�6$���ǅ �F��Z��4�
�X�B��M~rָm��.ة��y��D[�sc**I$���$C\��Z$?�1��e��Z@���Y%� ��a������H�V���5�럊^�C���j]��ь��Ge���\� '���<�\m�.�Tvark��h�����Z�~� v����4�|z����L���P��\L[$�]'�֜�խW���W�S�\Ҵ�U��)�IV�������۷Ƈ�6�}�rY���v�v�F7��+�~��
��B�O�5FG�'��X�^D�8��-R��-�F��V�A;uCl�V��sj,��'0s����5�>����X�
��
��� Y�Y�����! ��1��>��Y���>�Tp� �u���tt�v��K��F�p_%`W(o�=�Y��5X�-4���/&F՘���p������*C������ ( ^ܡ[%���g�u��~�V�jl�yKd}B�L]H�L{?�p��8p;Ip��臝_I8WG�����e8g�p��9��������50�x �7,FJ�*���d+c�g��~��� �k�°� ���> t	�#u�6��HS�p�r��!��<vuRP$��0��sHg#
�=B/�2 ���^v#�Nj���$������|	'!~��ځГ����½���x��B�~��O2��΀�w��I���f��@�2����q:Yb���#E}�87�_J�r�ݐ, $?��?�i� .Kj��B  ����DtVW�~���i|̍7�d�E�*���uo���-^s����-i�#����tu�&�&�P�9_]t>�.�����Z�a i�f�`6���a�d+�a5������wS�sI�R��*�8�t��刮�m�V�!�5�V����]h��Y�]�v��� �	�惯"��� �&2%��V��������(���*�f�Ƈ9=}�_���Y=��u�	x����v�0���?
��w��#�@����z�J�}9ե{9f�.|#"T����#���V����(x%.*�&���ɤg���?B�Wh>����u>�>	ժ>>��>�)s�s����:�U;���x���ec�!��(~�.</@.����=���@YD� ������`@@h����/t]���)a�x] ]]$�o~�w��y3��z��r}){)�%�Ip�H]Hb��V�8,
�'�D�a�@�f������8.���.u.	+�..�w.����*l�RE�����]�!�j1�Dj�n�A��Hn#A��ε-�h�
��i�,%�U���`%��ht'����}]d�4�B Q �3��3��Fa����Ј��v�PE���$9�'h�q�%�1%�J+&�J$J�J�T�%V���HI�$ԡI�$I�%���II�`I�� ��t#�V.�}Ǩ���b�V�#��a���Y�Kr�@U2'���	�E@�&"'b���g��l��"'����$�0�	
� [��C�CLh"�.��B	 �X��%	<�x,;��:��� ��^�&��*A�(2�W;
;��=;�Z����� 0�i` ��IV���dI��b���ǆv��� �x�� � �Ğ�h�v�!���z�&�?u����� ��.^�%���[�X�2J� ���<7���>au�@�99u��p�#���!�t�1�3�6�z9[8�]�Ϫm=���U�*[�kOD�C�Xr5��Xm����X�X����X;�6�)���XH��X�X����X,�X8� �XL�XZ]�l���X-�Jа�L���x��<A�<P? �[[�[ [��P�[P���YԸ�{� K���%=�5�A.�0G0G�Y�2[G�4��+5+\*+8+:Uz+<+>+�=@+�+A+�T+L%N��P+R�{+T+�+U+�"�+�V\��]+^]+`]�+b��+c:q�+;��S=6�>.?�:AxC�?QE"�'R�'' ��"X�4 ���D�91Q�m 99r�u�C��t���?����CUE�!>�.�P��S����� �XU
d?�A�K�[&������ �
[�Jx��J[y�"�Ι[[PmQ[ �yD�d&DeS�Z(-x 7�mʽ,���&;< i�=�QN< ����`���-�~�-~��#Y�,PV�~�D u@����K]�v��5��������V�RP9��+�� ?�� �  ������؊Ċ��*�N�y.�	w���˄��k�h��dl�����kE��^�4�4�y�4��;�2���#�2*�/��H��^B�q5�&�⫘��"����wRPD��E��� 6�KWW���QV�;i��UX����-x�V;���[�p_�u}��8�+�t�d �)ؖ�g�E�C�/��J
+<b�N ��+�;�r	w;�r0�Y�dv�Z���t�&�t;%�I�D���SE#~8~=/v�O�V $OV�1�bN���cC����
�Bб-$4��  e>\�%!:�����,Yz�,#,�х����
o&�w)AAD���,@���f�DءX]��U-�M9Sr^ i7�\D\�B�y���̋�K��~�B r��F�YO���Fw�`�`g����W� ��6#�����l<N�� ���]���t9-��F���M��y,���%Bh;v  �̀z�.t��B��+^o�ʢ���w����PC|KZE?�(g��(n��~�$�ɷo��.$��)(��WWV�]�E
P` !]�MU�u_U�`�0�	]W��f���3���,�EX
c��U%(� ��0�!<s�� ��6�+��` ur���ׁ�~����s��M��L2����6�&^TZT��:�zH6�XT��C��+��۴J(6 ���T��zX���+�xC�L; � ��3��6�T�`�T�ތc� ���pظ 6NTa�t���>Xa P����T� 5���`T��T%�6s�Y��W�.�y& �, ��W��3�6�̒Ws �M6����c��..�6��3% �= t,� � �T�t����u0 ��b���T��������tH���A� �����D�r
�6�t�@Ky羞W��$� 	� F3��X��}jn�tHS�Jpf 	l � ��sNoLp� � ��_t�>qC����Y�� " � ���+%�>�T���T�T ��;�s
OO���������� Et����� :���%{�>mB�����iT#���[�Y��+�� �;Ur@���3��  E�V3��B 2���2���7��U�����=,^ÏHU�B8�Tt)0`�, ��T A���3��u�GG��`>�T���ыѿp;�� �]�< t ��<	t�<to#z�kGN���\X<"t$< �\tB��3�A�g �Ӌ������u��91+�\1'�1�Ou1�10�����T�G��  ���+�ģ�T��� �6�?CC�6���f/V��62���ت�� f�w�y���3���ދ�b�^{'����\�l3��s�z"��.4/�*!�4�R4�4���4͏��o&U�qU�4���A IB�t���&�>$���E��E�@$�������>W�	� _ ����.�T��3 @�I��<;Ct�~ EE8��NQ�]9V0W+�V��W�;�g�@�t��@0����_b���W�	,���8���%��I��@�!_)��  ^Tr59XTs% P �ر��ً�+���Ë؜Xr8�$�H���.� 2���r�
3ys�PH�� X� �ș2��   â�T
�u#�>�Tr <"s r���< v��Uט��U�< ������WV�U+ �����D�t	+}�@ XtG��964Vs�m�23 �v�D�$���->��˹���;�üU'��K�G�L ���bu��d���D���~�gHubށ��M�����l`(��N1F��$U�N,Uu3y�u���u-�U�u��X���\� S��^��G ��K��Ҝ��eu6etP�<+|9>�y@?�?H����~W�^�pvs

	7Y��E�� t����S��!��\�8�����Q�P=6iw=9�̅��������V*vL����o��w�G��OM�����.l���@!���҉�A( ^�  �+��D$<t�uF'���,F�z~PC�����c�;@t���ķk�DkH0�d�w�3������X�ǧ��|����X�9��|�<�%X�X�����X���������<~z�:� "X  �|0u<F0l �3@+u�6��+�"��a �> ucc�@�	��-u�HF�d��R�V���Xfm��8 }�'�
�أ8.u�y#�F*�*�M<**
���V=F0 t2=N5=h =��l�!� .]7LLluF��|�M4��J����=ED
=�G=<	��X�� �-c = � v���.��4}��c��X���9�i�4�8�z>A��5��Q
����~XV>�8�a)���x�	�Q����\�!�����Xt'�g"�^ .t>���Ð�.	�}/�0	�k�����:
��Nރ�r�t"@Ak- �87�URA��A�A��G��/��p��*����ж��� 	 �ot��N�B2�GE %u���+�PV�������#;||�.��uY�|X�G tO)@��M�|�{�|���
A��{|
֥���|BH��tI
pIu��F뙐h��B�W�
�c���tu ���W��:�*m�(^���5���/,8��tL$N�r�RL�'6�XG��uN�}$��u�-F-\���G~D��L��#�1{�F�+���WzA����2t!W�w	�X+�ȉN�3�R0R��I���X� ���<a|�, FGL�}�����NBX���Xmu��زm>�`66�#u�#��y�d$�^�� �?t,?���u^�Ck95~�2*�F��@��6V�	���u	�=V(�eEN+�x�96�t���z�^��l4�F;�~��FqJu�H+�B�uW��y�C����o2>�����ҍ��;�gt�&Gu��*N��B�� xH�t4?��v�6�X
�����`�JV`
,H�ub�0��Ef�u$N*#�~���Oh��PI��Du/���Ox�9�7������S8���=@u�w.RJ�WBI���~B��K6���X�w88ɹ֗*�g۠ �?��gg�B���T'w^WG�P�Z�^��@Z}^���*ataԏu(hu=�h�!h
hH�G�p;��(�u93Mt~# �X�x �(V��aUFFu+~5���<�>����$�N���t2J�D�M�=�_	"���j �J&W�<'�{��(3�5*�]�=Ψ����Q>��>jLa����W�+u6%���Ð�0����R�L��������x�X �N�� �*u��?�F�h�H�����+�0|5909#��ua=s`(����� ^��0��F0�%h9~�	���C?���z�8DV�N��t
:u����+�^��(X;�Tr� 	�*�F�tH��~
3�ѹ�3BfK �
 uFVy(�,,��6G,�C$%�$�N��gn!���D
�=�F�������Tr=dzz�����}Ny�0��nq�F3n�o�Y���f��Z�T�
 -J�� =� vH��� \� =(s�� g<'�.+�  <
t;�t����# �avİ ��0DM������^_�U�E �R��PSQ��+���P��r��6Y[XU�sC$s	��:�&�?R�������+�T�'��u������Q�%?�9J�C
��B) �B�Y�U;�s=+�������:��t5�g�W�JV���)��s��h��$�9��L��V�� �ƀ�����6PV��؎�$�	 ���  � At�������s�w p�����tBH;�s����4�k����G�� t��L��H�f ���ƌڌ�;  �t&�XV��&�^��V=xt%3UHa�X�u�X�XG 0e���&�;�t���;�S�Ta�7뼠 wj ;�t$@@��'�^��M�����NN�4�]��G&��� G�Q� E�+�IAA��&�K;ZVv��` 8��r�r��#�+`o�� u��:Y�RQ�[W��d��G��  �+�J�U�XYZ�SP3�w�R�Br� �D��Z[tҌ��VW�X8�^T FHu�S r'�H0.�6�TH�;�:�D)V�:80 ^s0���v�sD� ��ڃ�������H�钉�T4'B�Ћ %N��9LtAu����?:r9�ӎ���hN9R�&L����	١�м�3�r\(����l�׋���:�n-u��#+���5�� ��I�����	��]�@��6�E��Zlǡ��3�;rW�h3j-p/����^���ܴ�WV�/ h}�(7;��[����2�9*���V �W� �j���}�� |L���\� ����r7\W��KU����!� �,�F�͋v�2�!l
<&p�q���3��`�DD�V􍗾'���p�}
�6U�^�]�q�6qp�E
r������ys18I�_�a�W���;F��EB��E�E�NW�-�0,��Mx*�\����W	����H����R��������������~y�1���u

��]_{������M���U�������VW�^@8�!{�S=K�K��G HT�����Q�׎��N} ^E=^N�_���O�W�
s����A��	���
O8t3��ǂz3zܿ("����i��6�6�9����X 
ݞc����� ���
u�y
�-��I����3g0�m�� ���0<9v'H�  �u�O���D��D;(�r�X�"E�@i=�k� !��W�Wu,�6�	�  4T7����y*��o�WÃ�u(|$�>jV�;@S�#� g��lV[�1�>�3�=-"�����7s
���opG�����Z��~��V  ύq�� .8tK�m�����I6N�tW��Ar(P�PR�� ��T�ԡ�vW= w1�R�q����K�V��Y�Ȁk��l< ? ��F]ZX�X�  ˣ�W��WUWVQS3��0�L�Kc�H��X[Y^_] ,���6�.�WSQpR2�P�P�=�J%���#Y[�G�.^
��R�ֽu,Ȉf
�9<�2����*���n�v	@��w�7���	$^t{."S��a�� N�������S��8˜fz�����!/�@�����w�|���a�{r;#wr�2vND�^[<�b35a_�:��Ea�ai�_3_+tV
\����� [֏�A��	����  � |��PP��� � 0 ��� ����<�	�t�� @���u����L��J(t�3����V� � �^����� �[��W�_skOu  ��Ӿ���}�=U��uǋ��&nInval�id partion ta  ble Error loadin�g operat
sys��tem Miss,� $�a�3^QR� pU���C� �p) `i�% ;�|+�� $���B���a���aL��� Ku���a+�*8� ];N{�~O� ]8��	���u��,��
<&�� u7<P�д���<�yy^����LG��8��� �a"T6��
,���
�����vЩ���m��m*��i�Vq�`z��~�s�?�i��~WЊ�� wx&FO��N �u�Ʋ ��.Ҽ8!�o7T�Y�.�� ��= �MS Run-  Time Library - C  opyright (c) 198 l8, Microsof :rp %4.0d�:%3%��'w	!FAT,16 	2t	 UNKNOWN v��̅t������ �����vH���g?��B	�."/ �\[]:|<>+=;,�Q%c-��2.2s
7.7`�
-11.s �-8.8s!�&$�  %1$�KФ�c8c�49���V
/PRIE�XTLOGQS0TATUS?MBR  l:\� �? �.?�1R�� ���{	(	 .�x�.�
R�7��s�IS&�&:sv[�#26S0 WU�!9� uC� @�r<��t7�u	���&�AtN�.'<=u.��C�sŬ��C�NWP��y�t�6`�H�</t6"t`GuT&�G2�.9f��s!���CC��2� �i�e�C`(@=\�2�h	CS'ƌ��sA4��,t�,4,
��	@6]�66 ]_[l.�=�	����;��P2���	.��.��K�Rt =�P��� �� X��X���UQH�rOs�o	� �!s� ����.�.�WY]�&�~ 	�E��E�3G��rJ&��P�+�.X��z&|��q:|	|&;xt&��Ձ�q� ���mm
����W�}>�&��ec�&�E`X<u
	UM �Z<u�P<t�{�<t�<���><u7�@81�/�]/+
u0
9P&�Gt�'�	t���{h0�� _�p�� S=(%PSRW7 ʦ��[�_Z[X�B� 0��a�.�>#u��I���� i�&@��� t
*�.�>�w����}X�PV.���2<:u�`dN �K�sFF��^&VR��(蔼�r-Y1.���Z^�  <�s<ar<<zw8$��4` SW�>̖8tPQR 0�e�»��� �8 �!ZY�].�E �CC,�&�_[�PB��-�m<+>Bm-�F���P3�3r �S�B�r92� p�������� r,��c4���	�	�����	Ճ� ŀAr��[� [D�k�����҃�&�r&�'����� Ft`)�F-�u&;Lr6g';T�.w<�(r:w �2H�||
|��Ɛ�	��u�� �b�=b$�6���	��@�nFR�DuBt�2�r2�22�r��EXr�Ü�u�Ýp� �<0r<9wb�,0uɃ�
�u�FF	����&URV8��#�#�Vt����#R!q�%t6
p�u\F�\&:F�ݙRFKyE$EFK�&E�@9@t&�G  t�N"���srO	O�D$�:tzj>�2�]SV� /3^���@���`�� r.�
�t�L�n��la%uY.�`<���}.�,��uG��
)
=�g�	'�Wu���#�? 'C
�'��ds��l[^HE����@��^ ��6l.�<�  t�RP� 8���!XZ��3ɝ�<���t��y<�0t��,�<-t&E" �)�r� ��
 ���(�r �F뽊���F����sì�"Q��q�9��t��	N��'�N�����SQ<t-�)^`2%&�} �^3�&�]��9�k�	CN&:���/Yj[6��0S��<[ �6<	t2<,t1u�D� F:��RD�rCMݚ�zKK K.�E��S 7�.!�;ݕ/u�P G.�G��2�r�0�+�X��N0@�VS���'PQR nWU3��޸ c`b��]_ZYXGC�Cm����
��
��:r:Dw�)h�� �[^V�����q� 碁��_�� 
�H#$AF�DOVer!�s!6 (C)�x�#��1-94�x�0censed��at;ialPr2tyke &/Al�Mse2rv5�W3�Ɏ�3��.��/�HE�>F/PN�T`^�DB��$�	y�@>\��Z%T��R11h f�}
���$�  �
 ��7�#3l$j@��Upn�  �.A Q�P rY_! ���H��PV��9�6v�xc�D�Z3� ������Dʫ��0=�j= s�����
Υ�B� ���WU���r����0�t���]���X�VS3�3�uļ�����%��tN8�W�[=' wZ0+Ã�2�7Y����������f��T�v��r0럜+u)RUQ��P��/<�Xu	�ظ?�ػ��Y\��]Z����b[^�/"yP2��qX_wG�����t=uP��!|�T���t�"��85����Dd+���&;�ك�	I���r
 `!u &}p�2�9G�|  `QUWR��zH��6Q��N�G& e &�rZ�N_�͐�
ZT]Y����S>`CA<"p5,5w s�Y����!2�6s�t��R r箼=a�����J��� s�U��HR �	GIu���Wp7PS���� ���u+�K��[�{I3�-OA�޴@��Z(UP�@�Z X� X�B�&�=u ����UQ`�����Ys��!�;��"]q�� ' � ��e` �ƀu~�>}�  � ��W�>v& �= �t&:r�:E  w�GG��_Ï�3�@���6����	v`���7�0RAe�t9�u 0�|
,u�6�A�"�	u����m����e�4�t!��%� &8%�8�e:�u S�s�BIu� NV���t3M�> ��u+�D0��7<<0��6�4��>G�.B4IOO� W+��
�_Ys����Q�ʊu۳u#�^��	���:3�Vh9iQ
m-8�D�|�L<��t^nBZ �RN  rHY_]^p
�dDr���'��0���X��`��C��@��� � ��
�C��E<-۱u� �-�� ] I�|�D	:�v�*���t
V�T|T�u�<0E�8Ls*� �ъ$����8���"�A��Uu�*
�Y#͐YB�
�t�
<��u�RU�G�l�c�ˬ�>9��rh"d<��]60uxPAx\�h�s�EPK2`Bt�GA��+�D]�-0 H�4 u$"`��u��C$!�N�u��T�u&&9�*��+C�}��,(��&U*��+*�*莆�����-R��   �4 \  G�` 	  p�o ,n   -� Incorrect	��v 0�
%1 al�aady instledbytesva��il� L�disk˄amec�Y0N /C%figur��9 hd3 f�"usCw��ith MS-�.4�9FDISK<=#��� ��P 3   �H  _  v "Canno���2In�d{wYk�|�Noji�	xeu�p��#nt���f�$zwritŸ,Th�mai<� bo{c�aog�YNOT6.e[�pd�3�d.�
$�3!���a^5Exn� Nd%1%�$���p �$Parh�!��!��WV�  ~�E
P��]�M�U 0�u_U�<�	]W��
��������ĉEX
^_�;l�D�)Dg�DP��N,X_P� 04<R>,
� �u3-˓3!13�! !!F@ �DGS�etupg��x)"�K))�l��b.|3��V~�"W79H�'>29b$,SOp^n�sW61�H6]C6te"�5�`��L��c���Dtve��W9� ac�Yt9��$3$Del�S?Y4�5isplayrB6inama��b1P���6Es(c to exi� A8A'Choosގ�f%��LllowS@:&1*56ha!NicuInt�E-�� ;)�"":�<FI>*20YWARONING!_꧿ԣ@B sD�--G1���rd�� unlX��a6hs}9D�7#EA�n�c�j
y�[<S4H> ]�S���P��[0M�6Pm���A`Y),Ӯ.��-Y2e�2-8&�(s)�?�I24 t�.ur>o � 	��� ���SDGyou���shS$f�tKx�87umRs$�izea�*Խ��@kI��� �(<Y>/<N>)� �.tA�?�g�A�xq�ox3xl8 Statx�� TypcVolc{�xel��Mr��("�9	Usagep_ޜIIHj޼��O#c<I��>	׵�:V+:�V�V.fTo�
�`space�7drr�(1
<d = �8576�K!)G5Q0GC>MLo0ER��M�^�]��N8NL��	O8��8�4T ��cgZ��(%)X��4d�Ic���.!
{ ���SI>
m� ��� �@��nt�D�sj��c�85�ueQ1� �	�C=� "X0300Q�arv#�I$��~{0���9�`��-̯�{�6���6o�:7��EE�`0341�l�0gK��63��6��7�(,7�����e�G�'�B��8

K�l�jߞ_�a�(�)Rk�޽�=í�.?�m
Bg �'�;AmA�d6[�n��n�bh���du��az���6��(W3�3UY�_tDU��C�-�]G�j�C�kG.j�C�kG/�ԟ13K4��KN-
��j��K�W9i�-BC<��O^ataR��dAdwwi��b&lost.l7P2vsWhB
� 2#d]�o&�R[..���<�2`��VI>��L{.�^GZ�]Q� �6�G��&N�
�� ���1�������a�1��?��A����xʮ׳�� 7�>AF�Y2s6 �++�P�i21r[�"'��.	%�[����C:n�{�>��/�*X����Miw��Ii�;��� �ka�}X@��sX-��zyxˢܐ�{T_?�5����`�`W��0�o�/6,�F���̲�NV02�� �eH0Z�F8e j��]�3����II>;
;�202 [(�:@�]�02�:���O45����2-2 O��@�a��t�>t�#b/�N�� N�._A-��)�.q$df��.�f0���^@響�>1�M�3�nowv��� �bI�Ins�/p�s,8e�.ttY�4A:J�����any %wh}ْ/&�.K��	|3�L֯/CMZI��D��CW{3R� +14�C�E"^?~>\���d����z�֭_�O�4e24�T\/,@ �l�r��sv$�Wd{]V�e<��{C�finr>J�ww�*�V.8�.D����be�Z@�j<��d�ic�X���(x�� ���xadp�Y��.��Err}���ڵ�8/wr﬇/�Inc0H�$v_;��."Can���awXh n���w5kǑ��d.~���_��߷9v���:palLex�t�Cs,�;r?�<�C_���������9Requ��evަ�sRso�t�q.��qZuv�$V���n�SH,(ly �m~`�&1R��gs[25�l�Y��>��uyb`{�]š,���� ��.<�Vc�IV%out�`� ��(�tv1eA��c��k jYs�sigPt��j[��dt�Ril�Xe�"}�Ͷ2����G>y��$���a�olX�PP�$�ц��1>gm��e�Tk�Yd7��$pA O��"n-�~��1mr:m�,�c�hbe=�+{w�c�c<y<G�ll�d�a zBoҡ�yr��T���@��!�1B>UnqB[�c�zC�J�O+3\� InvTid��ry,��ػ�!2Z�S���� �bqU��n0ؽg�g��H;l]d�doe<�xch�m��E;e�o��/cҞ��g�oX;�B.V�e��o֐G���#|Ng�C�x'WB>MsÉG�r%�e1��} Seh3I�>"H�C.MSG�</(��h�ƖHB���n!I% * Remo�	 PR�I  XENIX!�EXTT�PC/a HPF�NOVEbLLCP/M� �%�	�&���'�(5{���)��h���3!*�i+�=(-o�^��.�;/c{��A1�2�74_5��{6d�ϼ�87��g�
8F�3�,9t��gJ:$4;�3}�<�q=�����??A1��B�D@�� E:��{F�i�=�����G]��{��HZ������{I6c�JM����6K�����DL�M����3�%N`�=��O,�3o�P�=3]���QK��3 R0R<RDRLR �TR\RdRlRtR|R l /t@� L � �^T;C_FILE_INFO>�1 b� ����T.Cs��A	 #��Z[�+ �S	*���BIxI� ���U(nP�ull) +- #7� 4�tj�]	(e�tHaLP��
.5��R�S� �7ׁ��	*	p�x<<N�>>��gR6O
-�vck o*�gflow Tt3i��g�di.�vi'by I�3 	!9!��*eugh"%bp�n.ronm�<).� ��Y run-ti�&�� �KE2Exa�poqf�Tǥ�9'1lC�@#Y*�Q��c���
�J��rM� g�RB���`  �� ���   ��O����P�4 P����Ì�H��� �>���G�R��H������� H�+�s*+����H��ڋ��R ���¬��N�  ��F��$�<�u���� <�umm�t��2cx����3�)`c����i��  �t&��� �t�� ��[@���a��○>��6���-E������֋ ����.�/�@�� 0�ʨ��!��L�3P��!�fF��nup t���0�2A2�  1�9R9n8[878�7�6n6H=�;�@9@  @�?�?1?�>�>�>�>  >�=�=%WqVkr�����  �۴n���0�t����r�  r�r�
�����������������������  ��������������  ���������  �������~�z�  v�r�n�j�f�b�^�Z�  V�R�N�J�F�B�>�:�  6�2�.�*�&�"���  ���
�������` �������������  ��������������  ��������  ������B�>�:  �6�2�.�*�&�"��  ���`�r7s�씋7:;�   � 2� �   ��  �   r��  �R������Љ  ��"Win386 DSVXD Device  (Version 1.0)  	DSVXD_DDB                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            MZ�      � ��X�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          U�� �-��
�  RP�# P�����
P�Z���>�s)+�P�6�� P���� P��P� P�{��� �D�v�v�?���t	+�P�����v�v����>�?u���F� G�F� �F���F�P�F�P�����>� t�����F� ;�F���F�P�F�P����>� u�=���>� ug�>� u`� P��P� P����+�P�6� P����� P�F�P�X���F��P����F�<Yt<NuˊF��P���=N u	+�P�'����>� tF���t?� P��P� P�g��+�P�6� P�V��� P��P� P�D��� P��
��+�P��
����]�U��3��V�N�F�~ tI�^�7�</u�|?u�+�P�6� P����� P��P� P����+�P�6� P����� �+�^]�U�� �,WV�F� �z+�P�6� P���� P��P� P���� P�'
���~�t�� �^���v�0�����t*� �^���v�0�y���t� �^���v�0�����F��F9F�}9�v���v�4����P�>���t��>�?t�W��^���~�����r���t1�P��P���+�P�6�� P����� P��P� P����^_��]�U��0 �!
�F� �F���F�P�F�P�H����,@���F� �F���F�P�F�P�(���~� t,+�P�6�� P�f��� P��P� P�T��+�P�6��F��  �� +�P�6�� P�/��� P��P� P���+�P�6�� P���+�P��P� P����� P��P� P�����F�P�0���F� i��,@�FҍFމF֍F�P�F�P�F�P����~� ud+�P�6 � P����F�*�P�����F�*�P����+�P�6� P�z���F�*�P����F�*�P���� P��P� P�P����]�U�� ��F�P�Z���F�@����P�I ��]�U�� �+�P�6�� P���� P�F�P����F�P����uӍF�P��P���]�U���D�^�:t+��F���,@�Q�F� �F�J�F�P�F�P�S���~� t-+�P�6� P���� P��P� P���� P����F� �F�J�F�P�F�P����F�D�F�	��,@�F�F�P�F�P�����F� t-+�P�6
� P�'��� P��P� P���� P�����P��j�P����P��j�P�d���F�P�4����j��F����F��F� `�F�P�F�P�F�P�������8�j�t-+�P�6�� P���� P��P� P���� P�$��� ��]�U��3����^� t"��@@P� ���t� ��F@@P� ��+�]�U��3���>� t��  �D�>� t/+�P�6� P���� P��P� P�
��� P�����P��P�g���v��P�Z��]�U�� �DV�v�5���FP����F���P����F��~��~B�F�F�@= ~6�P��P�G��+�P�6� P���� P��P� P�m��� �{�F�  �c�F��~�}G�^�����^��v8 u� P��P����+�P�6�� P�(��� P��P� P���� �$�^��v�8 s�!��F��F�9F�}�F�  �+�^��]�U��B �K�"P�F�P������F��F�P� P�F�P����u.�F�P��P�^����,@���F� �F���F�P�F�P�2����]�U�� ��V��,@�}��P�P���F��F�  ��^��󊄮��~�F��F�9F�|��F� �F�v�F�P�F�P�����~� u�F� �F�v�F�P�F�P���+��� ^��]�U�� �f�~ u�v�����F�F�@�F�F�F�F��F�F��F�P�F�P�o��]�U�� �&�F�F���n��~�
s�F�0��F�7� P�F�P� P�����F$�F�<
s�F�0��F�7� P�F�P� P�e���]�U�� ��V�>��u-�F�D�F� �F�  �F�P�F�P�����F�t�� ����>� t,�F��F�P�F�P����~� u�6�>��� P����F�`�b �F�`�F�
�F�P�F�P�|���)P����F�b�>bu�6����� P�D���F�  ��^�F�v��F����F��a�9F�|�^� ^��]�U�� ���F� b�F�P�F�P����� �F�����&��F�<t	<"u� �+���]�U�� ��>� t�F� ;�F���F�P�F�P�����]�PQRSTUVW������+�P���_^][[ZYXϴ0�!<s� ���6 +��� r� ��ׁ�n�s��3�P�v��L�!���6�&26�&.�Ʊ��H6�,��6 ��+��۴J�!6�����p+�3���; ��3��6��6��6���P�� ���ظ 6�0tP�{���� P�0�0�!��� 5�!����� %���!�(�.��&�6, �*��3�6�&s�M6�.�ڻ 6�&��&�, �6��3�&�= t,� ���t��3��u������������tH���� ����� D�!r
�t���@Ky�2�2� �2�2� �U���R�} �2�4�t �U��4�4�f �4�4�l � �t�~ u�F� � � ���t�>�!C��� �F�L�!�(�� �&��� %�!�>� t�����%�!�;�s
OO��������;�s���Et����� U��� P�{�>� t���� P�i��]ø �[�Y��+�r
;�r����3��E�V3��B 2���2�����Ut��� P�,� ^Ï�� 8�t)��&�, ��3��� �3��u�GG�>������ыѿ �� ���< t�<	t�<to
�tkGN�< t�<	t�<t\
�tX<"t$<\tB��3�A�<\t�<"t��Ӌ���Ѩu��N�<t+
�t'<"t�<\tB��3�A�<\t�<"t��ۋ���Ѩu���>��G��׀��+�ģ����6�?CC�6���
�u��� 6���3���< t�<	t�<u� 
�u�y�6�?CCN�< t�<	t�<tb
�t^<"t'<\t���3�A�<\t�<"t�\��Ѱ\���s�"���N�<t.
�t*<"t�<\t���3�A�<\t�<"t�\��ٰ\���s��"���3���  �&�U��U��3ɋ����I�6, �t��&�>   t�E�u�E�@$������W�	 � _�ϋ���.���3�I��<;Ct�~ EE��
�u���N ]��]�U��VW�V�<�;�t@�t�3��������_^��]� U��W�v����t���3�������I� �@�!_��]� ��2r59,s% P�ر��ً�+���ËشJ�!Xr$�H�,��.22Ë���r3���]�s�P� X��]�s� ������]�2�� â�
�u#�>�r<"s< r���<v���ט��Ê���U���WV��+����D�tV�0��@tG��96s��^_��]�U���WV�v�~
�F�f�F��F��~ t�~ u+����Eue�߁���������������uL�F��u �v�V�E�P����F�=��t�+��v�� ��Mx������W��P� ���E u�F�N��Eu@�߁���������������t\�%�Mx������W��P�l ���E uSF�N��~� tI�} tϋE+F��#�F��F�PV�5��	���F��)F�)E���v�V�E�P�����F�=��t)F��F�+F��4��^_��]�U���WV�v�D��F���-�������������F��D�t�D@t�L ������Du�L�d�+��D���~��Du_�ށ���������������uF���t�� u3�v�����u-�����u�`���n�D��^��G ���V� ���Du�ށ���������������tP�<+|�D@��^��GH�D�~W�t�v������F����^���� t� P+�PPS�,���\�F���� ��P�FP�v�����F�9~�t����F*�^_��]ÐU���V�F-�������������F�� P����^�G�t�O�^��G ���^�O�F�@�G�^��G �^��D��G  ^��]�U���V�v�����u�F�`���� u$�F�n�Du�ށ���������������t+��5��-�������������F��F��D��^�� �G�D��L� ^��]�U���V�~ t[�~�t�~ uv�^�G�P����td�F-�������������F��v�K ���^�� �G  �^��+���G�*��^�`t�nu�G�P�[���t	�v� ��^��]�U���WV�v+��D$<uF�Du�ށ���������������t'�+D�F��~P�t�D�P� ��;F�t�L ����D��D  ��^_��]�U����^;�r� 	�*�F �tH�~
 t3ɋѸB�!rK�F
 uFVy(� ��6�V��F��ѸB�!FVy�N��V�� B�!�؋V�N�F
�B�!r������U����^;�r� 	��w���� t�B3ɋ��!r�����tn�V3��F��F��WV����f��N�T�
�uJ�� =� vH���ܺ =(s�� +�ԋ��N�<
t;�t����# �a�;�u� ��
�F���� ��^_�U�E3��e�PSQ��+���^�@�!rF��tY[X��Ã�s�	����@t�^�?u���� ��F�+F��f�^_���N�u�����V�@�!s�	���u����@t
�ڀ?u����� ��Y��;�s+�����3���U��^�t�O���]�U��VW�
�? u)� �su3���$@$��
��� ���D����6�N�؎��	 _^��]��� At�������s�w�����tBH;�s���t4� ���D����t��L�+�H����L��ƌڌ�;�t&���&�=��t%���t��H;�s����t�� ���D���G�t���&�t�،�;�t&��7뼋w3��j ;�t$@@��^ t�M�� t�NN뙌،�;�t&���G3���Q�E��t+�IAA��&;v��u����r�r��#�+�� u����u�3�Y�RQ� tW������D����w��+�J�U�XYZ�SP3�RRP� P� �����Z[t�� U��VW�~ u8�2�V�FHu�S r'�H�6�Ht;�t�D�FV�: ^s0�����s�u������ڃ��۱��H�!r钉�T�6�3�_^��]ËN��9Lt�����u���?��r9�ӎ�;�u9,s&����������;�u	١�+؎��J�!r;�u�,�����U��׋ތ؎��~3�����u��~������+����F�� t�I�������]� U��׋ދv���؎�3������ы~�Ǩt�I�������]�U��׌؎��~3�������I���]� U��^��!t��-  ���]�U��^;�}�� |���@t� �3���]� U���WV���v������V�b����F�VW� P�v�R����F�V�v������9~�u�Lx
�
����V�
 P�b���+������^_��]ÐU��VW�~��]�M�U�u�}
�!W�~��]�M�U�u�E
r3���u�� ��u_^��]� U��VW�~��]�M�U�u�u
�~��]_�!W�׎ߋ~��E�~��]�M�U�u�E
r3����� ��u_^��]� U��^�_��O�W��]� U��^�ӊ
�t,a<sA�C�
�u�]�U��׋ތ؎��v�~�ǋN��t�I�������]�U������U��3��ȋ"��Rt�"�F��t3���]�U��O�V�U��N�V��!��Nu�V�N���!�6�U��F�V�%�!3���]� U���!@� �^�3�]�             MS Run-Time Library - Copyright (c) 1988, Microsoft Corp  Incorrect DOS version
 Cannot label a JOINed, SUBSTed or ASSIGNed drive
 Invalid characters in volume label
  has no label Volume in drive   is  Volume label (11 characters, ENTER for none)?  Volume Serial Number is  - Delete current volume label (Y/N)?  Creates, changes, or deletes the volume label of a disk.
 LABEL [drive:][label]
 Cannot label a network drive Invalid drive specification Incorrect drive syntax -  Cannot make directory entry Unexpected End of File Multiple drive letters specified Too many characters in volume label
 Drive letter cannot be inside volume label *?/\|.,;:+=<>[]()&^"  ?:  ?:                              �      ??????????? m ��       CON �  �  ��       �  �  �    
 � @ �?:\ � B C [ � � � � � !E�����?e \      ?:\*.*       �  �L � L �2;C_FILE_INFO �  � ��� �  ���C �  �p   	��  `
  `
                   �      B � x �   � t �� �  �       � 	 �((((( �  �H � ��
 ������� � ������� � �  � � � �  �d<<NMSG>>  R6000
- stack overflow
  R6003
- integer divide by 0
 	 R6009
- not enough space for environment
 � 
 � run-time error   R6002
- floating point not loaded
  R6001
- null pointer assignment
 � �� ����������
    ^ �BRB��� �  ��� ��O����P�4 PˌÌ�H�؎�� � ���G����H��� ��������+�s��+�����ڋ������+�s��+�����¬��N���F��$�<�u���<�um�¨t��2� �3ҭ�����Î�������t&��� �t�� �܌�@����&H����Ë> �6
 � - �؎��  ��֋����.�/�@� � �ʎں�!��L�!Packed file is corrupt  �
D 	��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 MZ� @     ����    �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      U�� �K@�F�  �0%P��*P�k���<%$<u�0%PP�Q��� P�K?���K+���,��.�,,��,�v�v�(���F��t�62,P���� P�?���>�. t�9��.�# P�V����,��,��9�  RP�# P�V����*X�0%P��*P�T���t  �0%�F�
�u��*X��* �0%P��*P�T���t �X�F��~� u��*X��*  �0%P��*P�lT���t �6�,�6�,�# P�0V���~� u!��,,�t= t= t
����4,��!�v��4>��]�U�� ��>�F+ұ�=W�F��V��F�F��F�  �F�F�V���:X��]�U�� ��>V+����.��.��.��.��/�/� /�/��/�/�/�/��/�/�/�/�� /�"/��.��.�(/�
/�/��3�*/� :�:�$:�":�(:�&:�F��	 �n���ƇJ+ �F��~�|��v   �F�  � �n���Ǆ,/��+����4/��6/��0/��2/�v���晉��3���3���3���3����3���3���3���3�F��~�d|�^��]�U��
��=VƆ�� �F� �'�^���v�0����P�*P���~ P����P�P���F��F9F�|э���P��S�������2,�2,�? t1������P�� P�cS���t�2,�2,�����
�uڋ2,�? u+����?/tf��+��F���N��~� |
�v�����/u�F��}+��F���2,�2,�����
�t�P�� P��R���tދ2,� �v������2,� ��2,�G�-? = v�:��.����>,, t�2,�G � �Q�,, � P�� P�2,@P��O���uR�	 �P�>,, u��,, � P�� P�2,@P�O���u)� �'�>,, u��,, � P�� P�2,@P�sO���t1� 2,���>�. t�o���. � P�� P�2,@P�BO���uϸ �̓>�, t�C���, � P�� P�2,@P�O���u�� 롃>,, t���2,�F��,, � P�� P�2,@P��N���u� �� 2,������P�� P�Q���t�2,�2,�����
�u��F�  �(�����P�� P�[Q���u"�^��62,����,�2,�F��2,�����
�uʋ^�Ƈ�, �~� t����*m ��*��0%P��*P��*P�C���8%�F���*�F������F���^�������F��F��^�&�����
�u�^�� �����2,� �p�>,, t���>�. t����F�,�� P�v��	���F��~�2~�+�P�9���	��2,�G � �'��b�������������6���^��]�U��3��I:�FFu��*  �6�F�V�M(�O(�K(�L( �Q( �R(�S((�T(�U( ��* �F��*��* ��* ��*��*K(�0%P��*P� ��]Ð���Úp�Ú���3��9�d� �U�� �9V�(/���5�t+��/�/�/�/�3��* C��*P�0%P��*P�/ P�N���>0%�t� ��*C��*P�0%P��*P�/ P��M����*�F��2%�F��v�P�5����F��V��v��v���4����F��V�� �RP�v��v��P�:� �RP�v��v��P� :� �RP�v��v���O�":� �RP�v��v��P�$:��*R��*P�0%P��*P�*N����*��,�2%��,��,&�E u�H&�GE+ұ
��P�/�/�<%  ��* ��0%P��*P� P�0L���0%+ұ
�P��.��.�t�1+ұ
�P)�.�.��* ��0%P��*P� P��K���0%+ұ
�zP��.��.�J4�u� �G5�
�aP�/�/�2�u��� /�/)//��*3�0%P��*P�M���>7%u� �+����>7%u� �+���ƣ(/�|= ~
+��
/�/�$��*J�0%P��*P�/ P�JK���2%�/�
/  �>(/ u���P��3���t����+��(/�u��3^��]�3��S7�y 
�tt��* B��*P�0%P��*P�g P�K���6%+ұ�tO�/�/�2%+ұ�cO�/�/��* F��*P�0%P��*P�g P�K���0%*�%� ���&:�0%*�% �(:�U�� ��6��*5��*g��*P�0%P��*P�L���>�* t<�>2% t5�F�F��V�� P�v��
 P�6�*�NL��
� P�HP�F�P�I���t+��V��* @��*P�0%P��*P�g P��J���1%*�F���* F��*P�0%P��*P�g P�J���0%*�F��~� u�=@ r�� ��]�U�� �6�F�P�F�P��1���F��V��tQ�/�/�/�/�/ �/�F��V��F�V��%�^�&�?u&�G&�W�
�N//�N��F�
�~� uՋ�]ÐU�� �5V�F�  �F�F��F�F���F��^��?-u�N��F��^��?,u�N� �F��^�������O"t�
 �n��F��^���-0 F��׋^���F�<lt<Lu�N��F��^���F�<xt<Xu�N��F��^���F�<dt<Du�F��^���F�<ct<Cu�N��F��^���F�<st<Su�N��F��^���F�<mt<Mu�N��F��F�� �n���Ƅ@(ƄA( �F���F(�F���H(�F���I(�F�tJ�N��F��^��G���*��*��0%P��*P��*P����� �n���8%��B(�ށ�B(��*�GƄJ( �@�F�t� �n����F��^��G���B(��D(���F�� �n��؃F��v��D���B(��D(�F�t� �n���ƇG(�V�F�t)� �n���ƄJ(0�F�tƄG(3�6� �n���ƇG(#�'� �n���ƄJ( �F�tƄG(1�� �n���ƇG(!� �n�����G(�F�t*���� �F� t�@+��F��F�F��^��?%u����F��*��* �F���*��* ��*��t��*K(�0%P��*P�J����>|  u��|   ^��]�U�� ��2�^��W �� �
�VLRP�RP�F�P�G���^�Gu �v
�v�F�P�v�v�YP� P�����!�v
�v�F�P�v�v�v�mP�O P�������]�U�� �2�^��W �� �
��KRP��P�F�P�F���^�Gu �v
�v�F�P�v�v��P� P�����!�v
�v�F�P�v�v�v��P�O P������]�U�� �	2V��+�F��F�  �
 �RP�v�v��J0�^��F����$�
 �RP�FP�OJ�FFt�~�t�~�t�~�u�^��F��F����$�~ u�r�~ u��F�  �!�^����$�F��v�+�ƕ$����$�F���F��F��+���;F�ҋ^�Ƈ�$ ��$^��]�3��V1�>�. t9��.H��,;�,+��,  ��P�P P������D��P�
 P������,  ÐU��t�1+��F�F���*R��*P�0%P��*P�WF����*������,�2%��,ǆ��� Ğ��&��F+�H+  �>,,uF��P�
 P������P�T P������P�
 P�������P� P�������P� P������>,,uF��P�
 P�������P�= P������P�
 P������P�A P������P�B P������*0�0%P��*P�<E���>0%u�>1%(s�z ��z  +��F��F��F���F����RP�v��v�+�PP� P�����t� ��F�P� P�F�P�+ P�F�P� P��"���F�@ �F�  �F�� �F�  �� �RP�v��v�@ �RP� P����u��F�P� P�F�P�+ P�F�P� P�"���F�P �F�  �F���F�  ���RP�v��v�P �RP� P�E���t�S��F�P� P�F�P�+ P�F�P� P�/"���F�p �F�  ��,-p +ұ�=G- �� �F��V�RP�v��v�p �RP� P�����t����F�P� P�F�P� P�F�P� P��!����*  �>,,uY��,&�G"&�W$�
�^�&�&�W�F�V�=��t6��,;�s�R�v����P����P�A��� P����P��P� P����뵡�,�0,��,HH�.,�.,&��F��F�  ��,�F��F�  �v��v����+F�V���OF- �� �F��V�RP�v��v��v��v�� P�����t���F�P� P�F�P� P�F�P� P�� ���^�&�t��&�GF�@����ǆ��  S����F��V��^�&�G+ұ��E�F��V��^�&�St�� &�	Ct�� ��+�;H+|u;F+rm�F��V� �>,,t�1��P�
 P�����~�t��~� t���P�U P�w�����P�
 P�i�����P�R P�[�����P�S P�M������v��v��v��v��v��v�� P�����t����F�P� P�F�P� P�F�P� P����^�&�Hu:�v��v��v��v��v��v�+�P����t���F�P�0 P�F�P� P�F�P+�뵋F��V����������F��V����������F�P� P�F�P� P�F�P� P�K���F�@����ǆ��  �����9���r�Ğ��&�����<Dt<Iu
S�E�����P����P�>��Ğ��&��-B = w@��.����F�# �f�F�  �_�F�$ �X�F�( �Q�F�) �J�F�& �C�F�- �<�F�% �5�F�+ �.������������������������~�+u�<Ğ��&�G+ұ�C�F��V� �� �
�DRP��P����P�R?�����������F�V��^�&�G@F�Ğ��&�?Du3��@�F��F�  P�v��*��P��f�P�=���^�&�&�W�F�V��)���������"��P����P�f=����P��f�P�W=��Ğ��&�����<Dt<IuN�F��V�)�����������R�v��v��v���������� P�p���F�P�v��F�P+�P����P� P�b���>,,u$����P�v���f�P����P�F�P��P� P�w��Ğ��&�G@����F�9���v������������v��v���������� P������ �v��v������F��V��^�&�G+ұ� B�F��V��v��v�����P�>%P�R<���v��v�����P�~%P�;<���>%�^�&�G����ǆ��, �� &9Gu��@Ğ��&;t&�v��v��v��v��v��v��^�&�w�M���t�[��F�P�~%P�F�P�>%P�F�P�^�&�w����^�&�?Zu$�>,,us�u"��,P��P�G P�I���V�^�&�G@F�����P�I P�+���� �� �
�BRP��P����P��<������P�P��P�J P�����>,,uK�P�
 P������ �� �
��ARP�P����P�<������P�P�P�F P���� +���]�U��^ �'(V�P�
 P�����3�3u�P�Q P�j���?�P�a P�Y���P�
 P�K��� P�b P�=���!P�c P�/���F� �F�  ��F��V� �~� ~�� |	�~�dr�� �^���㋇�3��3u�� �^��㋇�3���3 �� �
��@RP�[���P�"P�F�P�;���^���㋇�3���3 �� �
�@RP�*���P�(P�F�P�c;���^���㋇�3���3 �� �
�z@RP����P�.P�F�P�2;���v����F�P���3P�F�P���3P�F�P���3P�F�P�4P�d P�+����^��]�U�� �&V�^&�G �t%�F�  �v��^&�@
�ވ��$�F��~�|���$ �U�^&�G
�= u��*A P�6j ��$P�:���%�^&�G
��*@ P��*A P�6l ��$P�p:���^&�G
��*��$^��]�U�� �&��*  ��* ���*P�0%P��*P� P�:���><% u6��*+ұ�5>;�.u&;�.u ��*�F��F�  �^�&����
�>�.�.��*b�0%P��*P��:���2%�F��F�  �0%P��*P� P�F9���0%+ұ
��=��.��.+��/�/�� //u	�//tX��.��. ////�F��V�+�� RP�v��v���<-  ���؃� �ډF��V���|�u�F��V��/�/��]�U�츒 ��$���t�� 9� t��
�t� �+��F��QP�
 P�2���RP�V P�$���SP�W P���+���F��V��F�V���.��.+�.�.�F��V�F�V���.��. �� �
��=RP�Z��P�TP�F�P�8���F��V� �� �
�=RP�2��P�XP�F�P�k8����.��. �� �
�=RP�	��P�\P��r�P�A8����r�P�F�P�F�P�[ P�`P�X P�R��� /�/+//�F��V�F�V�� /�/ �� �
�&=RP���P�oP�F�P��7���F��V� �� �
��<RP�}��P�sP�F�P�7���/�/ �� �
��<RP�T��P�wP��r�P�7����r�P�F�P�F�P�\ P�{P�X P����F�V��F��V��/�/�F��V�F�V� �� �
�t<RP�����P��P�F�P�,7���/�/ �� �
�K<RP�����P��P�F�P�7��+�PP����P��P��r�P��6����r�P�F�P�F�P�i P��P�X P�����/�/+//�F��V�F�V��/�/ �� �
��;RP�M���P��P�F�P�6���F��V� �� �
�;RP�%���P��P�F�P�^6���/�/ �� �
�};RP����P��P��r�P�46���~� t��r�P�F�P�F�P�p P�����r�P�F�P�F�P�] P��P�X P�)����P�W P����/�/�.�. ////�F�V�/�/�.�.//�F��V�F�V� �� �
��:RP�H��P��P�F�P�5���F�V� �� �
�:RP� ��P��P�F�P�Y5���F��V� �� �
�y:RP����P��P��r�P�05����r�P�F�P�F�P�_ P��P�X P�A����P�
 P�3����.��. //�F�V��.��.//�F��V�F�V� �� �
��9RP�x��P��P�F�P�4���F��V� �� �
��9RP�P��P��P�F�P�4���F��V� �� �
�9RP�(��P��P��r�P�`4����r�P�F�P�F�P�` P��P�X P�q���. /�"/ �P�
 P�Y����*n ��*��0%P��*P��*P����8%��n���*��p��//u�� �/�/ �� �
�9RP���P�P�F�P��3����p���n��6/�6/�k��P�P�F�P�3��
�F�P�F�P�P�l P����/�/ �� �
�8RP�,��P�P�F�P�e3����p���n��6/�6/���P�"P�F�P�@3��
�F�P�F�P�,P�~� t�q ��o P�O���4P�
 P�A���~� t*�5P�r P�-���6P�s P����7P�
 P���� /�"/ �� �
� 8RP���P�8P�F�P�2����p���n��6"/�6 /�Z��P�<P�F�P�2��
�F�P�F�P�FP�Y P����$/�&/ �� �
�7RP���P�NP�F�P�T2����p���n��6&/�6$/����P�RP�F�P�/2��
�F�P�F�P�\P�Z P�I���>�, tp�(/�|i= d�/�
/ �� �
�%7RP���P�dP�F�P��1����p���n��6
/�6/���P�hP�F�P�1��
�F�P�F�P�rP�t P�����(/=��t9=��t�t= t"�}P�: P�����zP�6 ��{P�5 ��|P�7 �܋�]�U�츔 �Ɔp� ���t�� 9� t�,�
�t� �+��F��~P�
 P�P���P�e P�B����P�
 P�4����P�f P�&����P�g P���+���F��V��F�V���.��.+�.�.�F��V�F�V���.P�F�P��.P�[ P��P�h P����� /�/+//�F��V�F�V��/P�F�P� /P�\ P��P�h P����F�V��F��V��/�/F�V�+��F��F��F�P�/PP�i P��P�h P�[���/�/+//�F��V�F�V��~� t�/P�F�P�/P�p P����/P�F�P�/P�] P��P�h P�����P�g P�����/�/�.�. ////�F�V�/�/�.�.//�F��V�F�P�F�P�F�P�_ P��P�h P����P�
 P�����.��. //�F�V��.��.//�F��V�F�P�F�P�F�P�` P�P�h P�C���-P�
 P�5�����
�u��>,,t���, �.P�
 P�����*P�0����*��*�>(  ��* S�>(��*��*�,��*P�0%P��*P�g P��.����, �>1%�u� ��* L�>(��*��*P�0%P��*P�g P��.���2%��l�ǆn�  �P��l�P�x2��p� u!�/P� P�r���0P� P�d��Ɔp��>�, u�1P��,P�,����l�P��,P�>(P�:P�, P�/��
�>(�>>( }�(��FP�
 P����//u�� �/�/ �� �
��2RP�t��P�GP�F�P�-���F�P�MP�F�P�-���|  �SP� P����F�P�/P�TP�l P����/�/ �� �
�2RP���P�^P�F�P�H-���F�P�dP�F�P�6-���|  �jP� P�R���F�P�/P�kP�~� t�q ��o P�1���~� t`�uP�
 P����|  �vP� P�	���wP�r P�����|  �xP� P�����yP�s P�����zP�
 P�����>,,u^��.��. �� �
�1RP�{P�F�P�r,���F�P��P�F�P�`,���|  ��P� P�|���F�P��.P��P� P�f���. /�"/ � /�"/ �� �
�K1RP��P�F�P�
,���F�P��P�F�P��+���|  ��P� P����F�P� /P��P�Y P�����$/�&/ �� �
��0RP��P�F�P�+���F�P��P�F�P�+���|  ��P� P����F�P�$/P��P�Z P����>�, tq�(/�|j= e�/�
/ �� �
�|0RP����P��P�F�P�4+���F�P��P�F�P�"+���|  ��P� P�>���F�P�/P��P�t P�(���|  ��P� P����(/=��t+=��t�u�� = u�� ��P�: ���P�6 P������>,,t�� +��F��F�9:tZ��P�
 P�����6 :�6:��P�F�P�u*���6$:�6":��P�F�P�_*���F�P�F�P��P� P�y����F� �F�  �>&: tT�F�F�u��P�
 P�R����6(:�6&:��P�F�P�*���F�P��P� P�*������P�5 �6���P�7 �,���]�U�� �V�F�4,�4, �6n �v��C(���^&�G�F��u�6r �v��)��� �~�u�6p ��F�H�F�F�V �F��V��F� �F�  �B+����~� }� �+��t'�~� t�F�  �~� tV�F�V �F��V��F�  �!�F��F��~�}��^�&��F�<u�� ��F��~�}�^��F��v��F�&����^�� �>z  t�v��v��v�� ���4,^��]�U�� �V�F�4,�>z  u� �0,9Fs�>4, t� �6r �4,P�(��� �F�F�F, �F��F�  �^�&�? u&� t�F���F��F��F��V��^�&�?uN�F���^��F��v��F�&���^�&�? u�^��F�� �~�4,v�^��?.u� �^���F�<\t<:u�F��v��4,P�&����N���^��]�U�� �V�F��'��' �F�� �^&�u�F�/ &� u�F�0 &�G�F��0,9F�s�~�� u9�F�+ �2�F��F��F�, ��@;F�u�F�1 ��F@�^�&;u�F�2 ��F�3 �F���*��*��0%P��*P��*P�Vك��8%�F���*�F��F�  ��^��F��v��F�&����'�^�&�? u�^��F�Ƈ�' �F�^��]�U��4 ��V�P�
 P�,݃��P�; P�݃��P�
 P�݃��P�? P�݃��P�@ P��܃��F�  �N� �Fָ �nԋ���0/��2/�4/�6/�FЉVҋ�0/��2/ �� �
�+RP�5���P�P�F�P�n&��� �nԋ؋�4/��6/ �� �
�+RP����P�P�F�P�<&���FЋV� �� �
�\+RP��߃�P�P�F�P�&���~� t,� �nԋ��F�P��4/P�F�P��0/P�F�P�F�P�vָ�f� �nԋ؃�,/u�	 �n�J+�� �nԋ؋�,/H�F��F�  P�v�������F� �nԋ��F�P��4/P�F�P��0/P�F�P�F�P�v�7P�N P�ۃ��Fԡ*/9F�}T� �nԋ؃�,/r� �nԋ���,/u��./�F�= t��F�  � �nԋ���,/t�o���4/�6/u�\��E �Y��F�  �� � �nԋ؃�,/ t�� � �nԋ���0/��2/�4/�6/�FЉVҋ�0/��2/ �� �
��)RP�TP�F�P�$��� �nԋ؋�4/��6/ �� �
��)RP�[P�F�P�$���FЋV� �� �
�)RP�bP�F�P�k$��� �nԋ��F�P��4/P�F�P��0/P�F�P�F�P�> P�iP�N P�eڃ��Fԡ*/9F�}��^��]�U�� ��V�~u��F��)�FH�F��F�  �6�S���F��}�F� ��F �F�V �>� t�~ u��������+�������  �� 9Fu5���t�F
Fu�������F  �� +������(�~ u�F
Fu�F�V���+�������F�  ��F��*/9F�}� �n����F9�,/u�= u	��./9F�u֡*/9F�u3=d u��P�D P�/ك�� ��� �n����F��,/�F���./�*/�>� t�F
Fu�F�V���F+�H+9Vv� r9Fr� � �n��؋F�V�0/�2/�~ u�F�V�.�.�~ u � /�"/9Vrw9Fv�F�V� /�"/�>� t"����9"/|9 /s�F�V� /�"/����9"/p|9 /sh����� /�"/�X�F�V //�~ u//� �n��؋F�V�4/�6/�~ u �$/�&/9Vrw9Fv�F�V�$/�&/�F
Fu+�� �v
���F�V��3��3�~ u0�F�V��3��3�F�V9��3wr9��3s�F�V���3���3�^
��㋇�3���3�F�V��t�F�V9V�r�w9F�v��^
���F�V���3���3�m�^��]�U��6 ���~t
�^
��W �>,,u�~t�v�v�v
�v�v�ك�
�>,,uc�^�GuY�~ t�� 9FuK�^
��W �� �
��%RP��P�F�P� ���F�P�v
�v��P�C P�փ�
�^
��W�>,,t��~u�6�F�P�����FʉF��V��)�F��*��*��0%P��*P��*P�(҃��8%�F���*�F��v��v������v���,P��!���t�0�uJ��P�
 P�փ���,P��P�< P�փ���P�
 P��Ճ���P�K P��Ճ���P�L P��Ճ��^
��W �� �
��$RP��P�F�P����^�GuF�~t�v�F�P�v
�v��P�H P�Ճ��m�v��v��v�F�P�v
�v��P�j P�hՃ��J�~t �v�F�P�v
�v�v��P�M P�BՃ��$�v��v��v�F�P�v
�v�v��P�k P�Ճ��^
��W�~t
�^
�/�_ ��]�U��( �
�^
��W �>,,u�v�v�v
�v�v��׃�
�>,,uc�^�GuY�~ t�� 9FuK�^
��W �� �
�#RP��P�F�P�W���F�P�v
�v� P�C P�oԃ�
�^
��W�>,,t�� �v�����,P�v�����t��,P�v�����t�� �uJ� P�
 P�ԃ���,P� P�< P��Ӄ�� P�
 P��Ӄ�� P�K P��Ӄ�� P�L P��Ӄ��^
��W �� �
��"RP� P�F�P����^�Gu�v�F�P�v
�v�! P�H P�Ӄ���v�F�P�v
�v�v�1 P�M P�kӃ��^
��W�^
�/�_ ��]�U�� ���  P�v�����ىF��N��t�^�&� ��]�U�� ��E P��$P�]���F�V�F��V��F��F��V��F��F� �F� �^&��=B tA=F t=L tw=S u� =X t��^�&� P�G P��$P�z����$�s�^�&�7�J ����,&�G?*�����u&�G?*�P�M ��&�G?*����P&�G?*�P�P P��$P�,�����,&�G!�@ P�V ��F� �^�&�7�^�&�7�Y �ˋ�]�U�� �V+��F96v ~�6�	 ��J+P����u��|� �96v u�6�	 ��J+P�3���v ��^��]�U�� �bV+��F96v ~�v�	 ��J+P�3���u�96v ~������^��]�     �           VDISK  V3.3                 �       VDISK3.3�  @  �     @UVW�5�!� � �H9�u�, &�E����&��t@�� - _^]�PQRSTUVW���������>t  t�F�X�F�  �F�P�F�P����6�,�6�,�# P�W��+�P���_^][[ZYXϐ�@ �ش �� ��<w� � ��$�82��!s���G,�ڊG�VW�U���3��� �� �h �=�!s�h $�=�!s
�z �=�!rP�g5�!� ��q �	 ��t3��U[� D�!rD� t>�� @t8�Ў؋չ +��F��D�!r ;�u�F���=-|� �� �� �D�!�3�P� >�!X��]�_^�U���3��F��
�/�u9�F� �F�
 ��u�F� �� ��u�F� �� ��u�F� �� �F� �� � �/�t�F� �F�  �F� � � �/<u2��؉^��܉^��F� � ��F�/�t���KSW3ۋ����/_[�u�F�  �F�  �F�  �F� �b���/���u��/�F� �F�  �F� �A���/<u<�t�F� �F�  �F� �"��F� �F�� �F� ���F�  �F�  �F�  �F��t� ��]�U�� �^��]�U�� �^]�U��V�	C�/<Cu$&�?
u&�G��v�&�G�v�&�G&�W�3���^]�3�P��X% �= �t3��U��3�����]�U��VW�>�  u� C�/<�u�C�/�� �� �� �� _^��]�U��VW2��� ��_^��]�U��VW��V�� 3�Ht��_^��]�U��VW��� 3�Ht��_^��]�U��VW��� 3�Ht��_^��]�U��VW��� 3�Ht��_^��]�U��VW��� 3�Ht��_^��]�U��VW��� 3�Ht��_^��]�U��VW��� 3��u��_^��]�U��VW��� 3��u��_^��]�U��VW��� ��º  u��_^��]�U��VW�	�V�� ��º  u��_^��]�U��VW�
�V�� 3�Ht��_^��]�U��VW��v�� 3�Ht��_^��]�U��VW��V�� �Kt��_^��]�U��VW��V�� 3�Ht��_^��]�U��VW��V�� ��º  u��_^��]�U��VW��V�� ����º  u��_^��]�U��VW��V�^�� 3�Ht��_^��]�U��VW��V�� �Kt���_^��]�U��VW��V�� 3�Ht��_^��]� �0�!�� � 5�!�� �� � %�vZ�!��#�.�� &�6, ��#��3�6��#s�M6��#�ڻ 6��#�� &�, �6��3�&�= t,� �� �t��3��u������ ������tH���� ��� �� D�!r
�t��� @Ky羺#��#� ��#��#� �U��$%�$%�} ��#��#�t �U�쾼#��#�f ��#��#�l � �t�~ u�F� � � ��� t�>�!C��� �F�L�!��#�� ��#�� � %�!�>�  t�� �� �%�!�;�s
OO��������;�s���Et����� U��� P�{�>�  t�� �� P�i��]ø �Y��+�r
;� r����3��V3��B 2���2�����Ut��� P�,� ^Ï� � 8� t)�� &�, �� 3��� �3��u�GG�>� �����ыѿ �� �� �< t�<	t�<to
�tkGN�< t�<	t�<t\
�tX<"t$<\tB��3�A�<\t�<"t��Ӌ���Ѩu��N�<t+
�t'<"t�<\tB��3�A�<\t�<"t��ۋ���Ѩu���>� �G��׀��+�ģ� ���6�?CC�6� ��
�u��� 6�� �3���< t�<	t�<u� 
�u�y�6�?CCN�< t�<	t�<tb
�t^<"t'<\t���3�A�<\t�<"t�\��Ѱ\���s�"���N�<t.
�t*<"t�<\t���3�A�<\t�<"t�\��ٰ\���s��"���3���  �&� U��U�� 3ɋ����I�6, �t��&�>   t�E�u�E�@$������W�	 � _�ϋ���.� ��3�I��<;Ct�~ EE��
�u���N ]��]�U��VW�V��#�;�t@�t�3��������_^��]� U��W�v����t���3�������I� �@�!_��]� ��Z#r59T#s% P�ر��ً� +���ËشJ�!Xr$�H�T#��.Z#Z#Ë��Qr3���]�s�P� X��]�s� ������]�2�� â� 
�u#�>� r<"s< r���<v��� ט�� Ê���U���WV�� +����D�tV����@tG��96"s��^_��]�U���WV�v�D��F���-� �����������!�F��D�t�D@t�L ������Du�L�d�+��D���~��Du_�ށ�� �������������!uF��!t��
!u3�v�����u-�� ��!u��%����,�D��^��G ���V� ���Du�ށ�� �������������!tP�<+|�D@��^��GH�D�~W�t�v��s
���F����^����  t� P+�PPS��	���\�F���� ��P�FP�v��6
���F�9~�t����F*�^_��]ÐU���V�F-� �����������!�F�� P�B���^�G�t�O�^��G ���^�O�F�@�G�^��G �^��D��G  ^��]�U���WV�v+��D$<uF�Du�ށ�� �������������!t'�+D�F��~P�t�D�P�c	��;F�t�L ����D��D  ��^_��]�U��d�w�WV�v�����%�F�%�F� %�%  �%  �|�<%t�X�% +��%�%�%�%�%�%�%��$�
%�"%  �|0u<F�"%0 �3�<+u�%�%  �"��< u�>% u�%���$�	�<-u��
%F��P�����u�V�%P�f�����>% }�
%�%�أ%�<.u#�%FV�%P�<�����>% }
�% �%��=F t2=N t5=h t =l u�% �>% u�<LuF�< u��% ���% ���% �ӊ�����=E t
=G t=X u	�%���� ����-c = v���.���H�%��%��%�i��%��$  �
 P����Q�� ���%�%�>% u	�% ���%  �%�% �>%u� +��%�F�9%t'�%�F��>
% t	�%  ���.%�%�}+��%�%� P�� ���: P�����~� t"�>
% t�F�- �%�}+��%���%  �.%� P� ����� �/�+�P���*��� ����������>% t��N��G�= t�=%u���+�PV�������< t�|��>% uY� %�G tO����MZHvG`H`H`HjHvGjHjHjHjH^G�G�GjHjHPHjHrGjHjHJH�>% t�>% u� %�G u��F뙐�%^_��]ÐU���WV�~
t�%�>%t�>%u�%��W�F��V��%�*�>% t�%��F��F�  ���%���F��V��%�>�$ t�F�F�t�F�+�� %�6%�>% u*�~� }$�~
u�-F�F��V��؃� �ډF��V��F� ��F�  �F���vW�v��v��
���>% t!W�	���%+ȉN����0F��I���N�%���t<a|�, FG�}� u�>% u�%%t�~� u� �+�P���^_��]ÐU���WV�~ t� �%�F��^��%� �>%u�%��W�F��V��%���%��F��F��^��%�>%u�F�F�u�"�	�~� u	�"�F��^��F��V��F�V�+�96%t�%���^��F�&�? tF;�~��F�^��F�&�? u�>%+��>
% uW���V�v��v��o���>
% tW���^_��]�U����%�F��~gt�~Gu��*��F��>% u�% �~� t�>% u�% �6%�6%�v�6%�v��>"��
�~� t�>�$ u�6%�@"���>�$ t�>% u�6%�D"���%� %  �%%t�v��F"���t� �+�P���]�U��V�>% u/� %�Ox�F�7��*���S�v����@u�%���%^]ÐU���WV�>% uI�v�~B��6 %�6"%�w���@u�%��N�~� %�Ox۠"%�?��*��܃>% u�F%^_��]�U���WV�v�>% uP��6 %�^&��P����@u�%�F��N�t� %�Ox��^&�� %�?��*��҃>% u�F%^_��]�U���
WV�6%+��F��F��>"%0u9%t9%t9%u�"%  �>%V�a���F�+�+~�>
% u�<-u�>"%0u��P�����N��>"%0t�~�>
% t�~ t�F��_ �> % t�F��j �>
% u&W�����~ t	�~� u�5 �> % t	�~� u�= �v�V������>
% t�"%  W�a���^_��]Ã>% t�+ ��  P����Ð�0 P������> %u�>% t�X ���x P�����ÐU���WV�v�F� �<*u�%�?�%F�H��<-u�F���F+��<0|5�<909>%u�<0u�"%0 �����������ȃ�0��F�<0|�<9~�F�����^�?��^_��]ÐU���V�""�N��F�< t
:u�� ��+�^��]ÐU����^;� r� 	�*�F �tH�~
 t3ɋѸB�!rK�F
 uFVy(� ��6�V��F��ѸB�!FVy�N��V�� B�!�؋V�N�F
�B�!r��� ���U����^;� r� 	������  t�B3ɋ��!r���� �tn�V3��F��F��WV����f��N�T�
�uJ�� =� vH���ܺ =(s�� +�ԋ��N�<
t;�t����# �a�;�u� ��
�F���� ��^_�U�E3��
PSQ��+���^�@�!rF��tY[X��Ã�s�	���� @t�^�?u���� ��F�+F��f�^_�'�N�u����V�@�!s�	���u���� @t
�ڀ?u����� ��Y�� ;�s+�����3���U��^�t�O���]�U��VW�("�? u)� �su3���$@$��("�*"�� ���D����6."�N�؎��	 _^��]��� At�������s�w�����tBH;�s���t4� ���D����t��L�+�H����L��ƌڌ�;�t&�6"��&�<"=��t%���t��H;�s����t�� ���D���G�t���&�<"t�،�;�t&�2"�7뼋w3��j ;�t$@@��^ t�M�� t�NN뙌،�;�t&�6"��G3���Q�E��t+�IAA��&;8"v��u����r�r��#�+�� u����u�3�Y�RQ� tW������D����w��+�J�U�XYZ�SP3�RRP� P� �����Z[t�� U��VW�~ u8�Z#�V�FHu�S r'�H�6�#Ht;�t�D�FV�: ^s0�����#s�u������ڃ��۱��H�!r钉�T�6�#3�_^��]ËN��9Lt�����#u���?��r9�ӎ�;�u9T#s&����������;�u	١� +؎��J�!r;�u�T#�����U��׋ތ؎��~3�����u��~������+����F�� t�I�������]� U��׋ދv���؎�3������ы~�Ǩt�I�������]�U��׋ތ؎��v�~3�������+��t������]� U��׌؎��~3�������I���]� U��WV�N�&�ً~��3����ˋ��v�D�3�:E�wtII�ы�^_��]�U��VW� �U��^;� }�� |��� @t� �3���]� ����P#
�u�P#�����!� � U��VW��
�F�͋F�F�<%t
<&t�F����F���F�D�F�D�V�F��F�~��]�M�U�u�}
U�^�]�W�~��]�M�U�u�E
r3����� ��u��
_^��]�U���WV�F���F�F��EB�F�E��E��FP�vW������Mx*������W+�P������^_��]�U��VW��
�F�͋F�F�<%t
<&t�F����F���F�D�F�D�V�F�F��~��]�M�U�u�u
�~
��]_U�^�]�W�~
��E�~��]�M�U�u�E
r3����� ��u��
_^��]�U��VW�~��]�M�U�u�}
�!W�~��]�M�U�u�E
r3���� ��u_^��]� U��VW�~��]�M�U�u�u
�~��]_�!W�׎ߋ~��E�~��]�M�U�u�E
r3���3� ��u_^��]� U��VW�^�v�F�~
�N�_^��]�U��^�_��O�W��]� U��W�~��3�����A�يF���O8t3���_��]�U��֋v�^��
�t,��'C:�t�,A<ɀ� �A��,A<ɀ� �A:�t������]�U��^�ӊ
�t,a<sA�C�
�u�]ËN
�F�V�~W��
�t��
u�y
�-��ۃ� �ڋ��3��t�����0<9v'����u�O���D��D;�r�X_^��]� U��F�5�!�Ë�]�U��F�V�%�!3���]� U��WVS3��F�}G�V����  �F�V�F
�}G�V����  �F
�V�u�N�F3���؋F����8�؋N�V�F���������u�����f
��F���r;Vwr;FvN3ҖOu���؃� [^_��]� U��SW3��F�}G�V����  �F�V�F
�}�V����  �F
�V�u�N�F3���F���3�OyC�H�؋N�V�F���������u�����f
��f�r;Vwr;Fv+FV
+FVOy���؃� _[��]� 2��������� U��^��W�N����^��W��]�  U��^�v�v�w�7� �^�W���]� U��SV�F
�u�N�F3���؋F����8�ȋ^�V�F���������u�����f
��F���r;Vwr;FvN3Җ^[��]�  U��S�F
�u�N�F3���F���3��E�ȋ^�V�F���������u�����f
��f�r;Vwr;Fv+FV
+FV���؃� [��]� 2��������� �0�!<s� ���6 +��� r� ��ׁ�.:�s�;�3�P���L�!����6�&Z#6�&V#�Ʊ��H6�T#�6 6�R#��6 ��+��۴J�!6�� ���$�0:+�3���u�����;�3��6� �6� �6� 螥P�� �X#�?P���=�� P�X#          MS Run-Time Library - Copyright (c) 1988, Microsoft Corp %c: %c: - %c: ---------- IO     MSDOS   B F P [ b            	  /	 CLASSIFY DEBUG FREE PAGE ALL MODULE  :	  /	              ����        ����        ��������        ����       
     
 $A �MS DOS Version 6 (C)Copyright 1981-1994 Microsoft Corp Licensed Material - Property of Microsoft All rights reserved PSRW3Ɏ�3��.� �/�� �>� �.��/�� �>� �.��/�� �>� �.��/�� �>� �E��� �>� �� �>� �f��� �>� �.��/�� �>� �� 
�<$��   �� 
 �Y��� �>� � ��� �>� � �. �A Q�P rY_Z[X�����PV� c�!r�6� �� ^Xø D�  3��!�����D�!ø D� 3��!���D�!ô0�!=u��= s����� � �  � ����PWU���r����t���]_X�VS3�3ɀ��uļ� ���%��tļ� ���= r=' wļ� ���ļ� �Ã��u���u���� ���� 3����� t�T ���r�u럜��u)RUQWP� �/<�Xu	�ظ�/��s_Y���� ]Z�����[^�WP���2����IX_Ã�u�>� �t=��uP�� �� X��� �3ɀ��t&�M�	&85u&�M���s+��t���t&;�&;u�	It�����r
����u &}r2�&�G��  �PSQUWR��� �6� ����t�u�& ��rZ�_�����_Z�r]Y[X�����PSR�� ���u�, ��w s�Y�  �!2�������t;�t� ���rZ[X���u�&��!��� s&�U�!����t	&��!GIu���WPS���ٰ��u+�K��[X_�3��tO�@�׃�u(�!P&��Z Xs��@B�!�&�=u��������UQ����Y�!s�;�t;��u��]ø' � �À��t�ƀu�>� � � ��W�>� �t&�= �t&:r&:Ew�GG��_Ï� 3ۓ��6� ��6� ��	v��7���0RA�u�t9��u�|
,u�6A�"��u�|
,u�6A���u�|
,u�6A�3��3�3��6� �3��t!�%� &8%u
&8et:�u&��S�sGGBIu�V���t3M�>�  u+�D0&:Eu�<0u�t4��>� �uBBIIOO����W+��
�_Ys��Q�ʀ| t�tIIGG�^��u^�	���u3��tVUWQ3Ƀ>�  u-�Du�|�L��Dt�Dt�Du�|�Z� �R ��  rY_]^���
��>�  ur����   �3ҡ� �� 
 ��X��� C��@u�� ��u�
��� CC�� �3ۀ| uǇ�  -CCƇ�  C� ]3�3҈� �D	:�v*����D�t�D
��� C��@u�| ��u�| t8Ls*L�ъL�t$�Du�Dt&�G�X��� C��@u�A ��u��D�u
�t�D
��� C��@u�# ��u��Du�Dt�
�t�� ��u�� U�QW��3ۍ>� ��r_Y�����]�D0u&�PA�h�s&�EP��&�
�tGA��+�U�]3�3���  3��D u$&��Du��tC$�� 
 �Du�� 
 �T�Du&&��Du�ĀtC���� 
 �Du�� 
 �(&�&�U�Du�ƀtC���� 
 �Du�� 
 �D@t)PR�82��� �!s�,�D
��ZX�D
,����ǈD
�����t3Ҳ-RU��d �
 � � �  3 U t � � � �   # 7 E Y m m p y �  �! �" �# �$ �% �& �' �( �- �8 �9 �; �< �= > ,? .@ mA �B �C �D �E 'F +G <H YI qJ �K �L �M �N O /P MQ iR �S �T �U 	V W GX sY �Z �[ �\ �] �^ �_ �` a b  c Ud �e �f �g �h  	i 1	j 7	k Q	l j	m �	n �	o �	p �	q �	r �	s 8
t o
,�
-�
./�0R1�2�Incorrect DOS version

8  Segment^	�  �Total �  �Name � 	 �Type
<  ------- � 
 �- �   �- �   �- �
%  Handle      EMS Name      Size   
%  -------     7 �- �     ------  
"   %1 �  �%2 %3  %4     %5
' �  �%1 %2     %3  %4%5
0 � ( �%1  %2
+Memory accessible using Int 15h     %1 %2
  %  XMS version %1; driver version %2
  EMS version %1
	LOADHIGH Temporarily Restricted Interrupt Vector ROM Communication Area DOS Communication Area IO MSDOS System Data System Program System Device Driver Installed Device= %1: 
%1: - %2: 	BUFFERS= FILES= FCBS= STACKS= DEVICE= IFS= 	INSTALL= IBMBIO IBMDOS "Modules using memory below 1 MB:
#%1 is using the following memory:
Free Conventional Memory:
Free B  Name��  �Total       =   Conventional   +   Upper Memory
D  4 �- �   �- �    �- �    �- �
  Segment � 	 �Total
  -------    �- �
   %1    %2 %3
=Too much of memory fragmentation; MEM cannot work properly.
SYSTEM   Total Free:%1 %2
 %1 is not currently in memory.
   %1� �  �%2 %3  %4
% �  �- �
  Total Size:      %1 %2
+  Segment  Region       Total; �  �Type
/  -------  ------   �- �   �- �
   %1     %2   %3 %4  %5
  %1  %2 %3   %4 %5   %6 %7
!   %1     %2   %3 %4  %5     %6
Press any key to continue . . .No upper memory available
8  Segment  Region       Total� �  �Name � 	 �Type
<  -------  ------   �- �   �- �   �- �
Conventional Memory Detail:
Upper Memory Detail:
.Memory TypeC �  �Total  =   Used  +   Free
/ �- �  -------   -------   -------
%1  %2   %3   %4
+Largest executable program size     %1 %2
+Largest free upper memory block     %1 %2
Conventional Upper Extended (XMS) Expanded (EMS) Total memory Total under 1 MB Free Upper Memory:
8  Region   Largest Free     Total Free      Total Size
:  ------  8�- �   �- �   �- �
    %1   %2 %3  %4 %5  %6 %7
Memory Summary:
7  Type of Memory       Total   =    Used    +    Free
:  n �- �   �-
 �    �-
 �    �-
 �
  %1  %2   %3   %4
	Reserved    %1' �  �%2 %3  %4%5
   %1     %2   %3 %4  %5%6
+Total Expanded (EMS)? �  �%1 %2
module name bytes +Free Expanded (EMS)/ �  �%1 %2
Extended (XMS)* +Free Expanded (EMS)*- �  �%1 %2
@* EMM386 is using XMS memory to simulate EMS memory as needed.
:  Free EMS memory may change as free XMS memory changes.
+Available space in High Memory Area %1 %2
?Displays the amount of used and free memory in your system.

AMEM [/CLASSIFY | /DEBUG | /FREE | /MODULE modulename] [/PAGE]

�  /CLASSIFY or /C  Classifies programs by memory usage. Lists the size of
}�  �programs, provides a summary of memory in use, and lists
: �  �largest memory block available.
{  /DEBUG or /D     Displays status of all modules in memory, internal drivers,
r �  �and other information.
�  /FREE or /F      Displays information about the amount of free memory left
g �  �in both conventional and upper memory.
�  /MODULE or /M    Displays a detailed listing of a module's memory use.
s �  �This option must be followed by the name of a module,
7 �  �optionally separated from /M by a colon.
@  /PAGE or /P      Pauses after each screenful of information.
�>���}��) D * L + T , S . f / � 0 � 1 � 2 � 3 � 4 � 5 � 6 � 7 : A> u�wLASTDRIVE= � �-
 �       %1     %2     %3
/%1 bytes available contiguous extended memory
System Stacks -- Free -- Program Environment Data %1 bytes available XMS memory
$The high memory area is available.
(The high memory area is not available.
-MS-DOS is resident in the high memory area.
7MS-DOS is resident in ROM using the high memory area.
Free  �>d������ Extended Error %1�>+�� ��� Parse Error %1�>O���U��WV�~�E
P��]�M�U�u_U���]W�~
��]�M�U�u��ĉEX�E
^_��]�U��WV�~�E
P��]�M�U�u_U�!�]W�~
��]�M�U�u��ĉEX�E
^_��]�U��WV�~�E
P��]�M�U�u_U���]W�~
P��]X_W�~��]�M�U�u��ĉEX�E
^_��]�EMMXXXX0  (%ldK) %5lx%,8ld%7c%-8m%-m %5lx%3ld%,8ld%7c%-8m%-m (%ldK) %5lx%,8ld%7c%-8c%-c %5lx%3ld%,8ld%7c%-8c%-c��  �%-8c%-m        (%ldK)   %,8ld%7c%-8c%-m%-c %-c  (%ldK) %,8ld%7c  (%ldK) %,8ld%7cP �  �(%sK) (%sK) (%sK) %3ld%,7ld%6c%,7ld%6c%,7ld%6c    %sK %sK %sK %-16m%7c%7c%7c %sK %sK %sK %-16m%7c%7c%7c %sK %sK %sK %-16m%7c%7c%7c %sK %sK %sK %-16m%7c%7c%7c %-16m%7c%7c%7c  %sK %sK %sK %-16m%7c%7c%7c  %sK %sK %sK %-16m%7c%7c%7c  %sK (%s %s)   %6c%17c %sK (%s %s)   %6c%17c     %sK (%s %s)   %6s%17c %sK (%s %s)   %6c%17c %sK (%s %s)   %6c%17cW� 
 �%-16m%,10ld%,10ld%,10ld %-16m%,10ld%,10ld%,10ld %-16m%,10ld%,10ld%,10ld %-16m%,10ld%,10ld%,10ld %-16m%,10ld%,10ld%,10ld  %-16m%,10ld%,10ld%,10ld  %-16m%,10ld%,10ld%,10ld     � �  � %,5d%8c%6lx  (%sK) %8.8s  %,10ld%8c (%sK) %8.8s  %,10ld%8c       (%ldK) %8.8s  %,10ld%8c (%ldK) %8.8s  %,10ld%8c (%ldK) %8.8s  %,10ld%8c (%sK) %8.8s  %,10d%8c       %d.%02d %d.%02d %5c%5c  %d.%02d %5c      (%sK) (%sK) (%sK) %-8m%,8ld%7c%,8ld%7c%,8ld%7c %-8c%,8ld%7c%,8ld%7c%,8ld%7c (%ldK) (%ldK) (%ldK) %-8m%,8ld%7c%,8ld%7c%,8ld%7cL�  �(%ldK) %5lx%8ld%7c  %-c    (%ldK) %5lx%8ld%7c%-m %5lx%8ld%7c%-m%-c %5lx%3ld%8ld%7c%-m %5lx%3ld%8ld%7c%-m%-c (%ldK) %5lx%,9ld%7c  %-c    (%ldK) %5lx%,8ld%7c%-c %5lx%3ld%,8ld%7c%-c ? %d %d %d %d,%d %c %d,%d  EMMXXXX0EMMXXXX0 MICROSOFTEMMQXXX0� �  ��<  ;C_FILE_INFO �  � ��� �  �� �C �  �0;   	��  �(  �(                   �      B � x �   � t ��!(null) (null) +- # �  �     ^@^@^@^@^@        � 	 �((((( �  �H � ��
 ������� � ������� � �  � � ���      �?  � � L �Z# �  ��C<<NMSG>>  R6000
- stack overflow
  R6003
- integer divide by 0
 	 R6009
- not enough space for environment
 � 
 � run-time error   R6002
- floating point not loaded
  R6001
- null pointer assignment
 � �� ���������Y    v L	�RB��� �  ��� ��O����P�4 PˌÌ�H�؎�� � ���G����H��� ��������+�s��+�����ڋ������+�s��+�����¬��N���F��$�<�u���<�um�¨t��2� �3ҭ�����Î�������t&��� �t�� �܌�@����&H����Ë> �6
 � - �؎��  ��֋����.�/�@� � �ʎں�!��L�!Packed file is corrupt � �\�\�\�\t]�^ucu�u����9{b{�}�Y                                                                                                                                                                                                                                                                                                        MZ� *     v ��w�    �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      . .. 
 �JJJJJ����.;;;;;;;;;;;;;<;<�����������������;�CDROM CD001 $+: \NEWELL.DAN \.  ~ �  �  � �  �  �  ��           �  �EMMXXXX0 �  �� � ' �Zp����RS5S]S�S�S�S�S	T"T?TPTiT�T�T�T
UU/UDU[U�U�U�UCDR100: Unknown error CDR101: Not ready CDR102: EMS memory no longer valid CDR103: CDROM not High Sierra or ISO-9660 format CDR104: Door open� � �DN0:\DN  �� �  �<   G   �  �  �  �  �  �  �  �  �        $  6  :  J  P  `  �       �    _ �  �       �� �  ����DNMSCDEX  �  ���6 � ��U��WV�v�~��< tF��O�u�� ^_]� U��~ tD�^&�? u�  �F�^
�F �+�^&�?u"� �F�^
�F ��^�F&��^�F&��F�N�u��^&� ]� U����F�  ��F��^�F&�? u�F���]� U����^�F&��^�F&��^&�? u�&��^&�]� U����^�F&��^
�F
&��F�N�u�]�
 U����f�V�n�~ u�F�V]� U����n�^�n�~ u�F�V]� U����F�  �F+�;Vwr;Fs�F+�)FV�F��ߋF���]� U�����~�ar�~�zw�^&�/ �F�^&��F�
�u݋�]� U����^�_��� �F�= s= u� �� #F�f��+���]� U����^�_��� �F�= u�F�V��v�v� ��v�P����]� U��VWP���*X�v�^�\�v�\P���*X_^��]� U��V�v+��D��D�D�L�d��D^]� U���V�6 ��F9DuV������ �&  ;�u�^��]� U����^�Gu� �N�^�G*�F��F�t+���F�t� ��F�t� �� �F��^�
��� �G�w�v��q+�t�+���]� U���V�v�t�t�t
� P�v�v�[)�F��t+����F�V��T�F�^��]� U���
WV+��F�	 �6 �5�Dt���FtX�F�  �F�+F��F��|
u�D9Ev���F��F���� �&  ;�t"�Du�D*�F��F�"F�t��F9Du����u+��K+��E��
 �
 �E�>
  u�6 ��D  ��� �&  ;�u�F�E�e��F�EW����^_��]� U���V�6 ���� �&  ;�t�F9Du��T9Fu�9Vu�V�G����+�^��]� U����v
�v�v���F��t�F��&�v
�v���F��u+���v��v�v�d��t����]� �U���V��,�F9Du!�~ t�F9Du+��D�D�D��D
�D�����r�^��]� U���V�V�F�F��V��������s.�F��V�9Du�9Tu�������� ��T�D�T
�+��^��]� U���V��F����F����&��T9V�rw9F�r�v���T�F��V��t	�����rԋ^��F�V�G�W
�������� ��W�V�F
�G�W^��]� U����p�F���F�%�% �&np;F�t�^��F�V9Gu�9Wuً��+���]� U����p�F���F�%�% �&np;F�t�^��F8Gu���+���]� ��RP�z���F&�w&�7�k��U���
���J&��F��V�RP���u+��F�^�&�G,@�F�&�G,A�F��p�F���F�%�% �&np;F�tˋ^��F�8Gu�F�8G$uًË�]�U���^&���u&�w	&�w����+�]� ��RP�����B&�w&�7����+��U����*�F�= u+�
��F��V��^�&�:u&� ,`*�P����F��u+���]�U����"&�&��F��F�@t�F� t�6&�? u+���"&�&�$*�P�z���]Ë�RP�-��+��U����� *�F����㋇ �F��t�V��� �F�= w�F��=�v��~�t�~�t�~�t�~�t�~�.t�~�-u� �+�P���t��F���뾋�]�U���^&�G�^&�G�^�G"t�^&�G&�W�
�^&�&�W�^&�&�W�^�G"t	�^&�G��^&�G�^&�G�Ì� RP�F�V RP�^�G"t�^&���^&�G*�P+�P��]�
 U����~ t	�^&�G��^&�G�t6�~ t	�Ì�X �	�F�V` �F��V��x PR�v�� P�� �u� �+���]� U���WV�^�w�G"*�% �F��F� �F�  �v� P���F��t� +���~� t�^�&���^�&�G�F��~� t&�G��^�&�G�F��~��u�~� t��F�  뜀~�u;�~� u�~�u�~� u�� �^�O"�� �~� t�~�u�v��v��v�����u��v��v��v�F��V� �-��t�^��^�G
�W�F�V��r P�F�@RP� P��= ��ىN�l P�F�V�	 RP� P��= ��ىN��~� t���t�	��v�,�+�P�^�G*�P�`�� P�^�G��*�P�P= t������^�g"��F���~� t�^�&�GP&�WR��^�&�GX&�WZ��� ��� �~� t&�Gx��^�&��� ��� �~� t&�G|��^�&��� ��� �~� t&��� ��^�&��� ��� �~� t&��� &��� ��^�&��� &��� ��� ��� �~� t�% ��  �F��DP�~� t�F�V�( �	�F�V�0 RP�v����D'P�~� t�F�V���	�F�V��RP�v��}��DMP�~� t�F�V���	�F�V��RP�v��V��DP�v��u�D'P�v��k�DMP�v��a�~� t"�DsP�F�V�RP�v����DsP�v��;���Ds �F�  �J� ;F�~M�~� t�~������^�&��� &��� ��~������^�&��� &��� �^����㉀� ��� �F��~� t�� ��v�~� t�^�&��� &��� ��^�&��� &��� RP� P���P�~� t�^�&��� *�+�&�� &�� ��^�&��� *�+�&�� &�� RP�i �v��� ��� ��� RP� P�q�P��� ��� �C � ^_��]� U���>V�^�_��� ��� �FĉVƋ^�_��� ��� �F��V��vRP���F��V��v�v��v���F�+�F�VƉF։V�- �� RP� P���@�F�F��V�F�V�F��V��F�+ҹ' ��@�F��F�  �F�  ��^̀O�Fԉ�ÉF��FڋF�9F�s�v� P���F��u�+����^�F̉GS�v��v��F��V� � P���F��t��F� �^�G�F��r�^܋F�&�G&�G��+�&�G&�G�F�&��F�&�G
�F�+�F�V�;V�r?w;F�v8�^̀O�v�v��v��F��V� � P�2��F��u�]��v��\�^̀g���F�  �^̋G
�WF��F�V��G
�N֋^��u�� v+۹ ��F�V��F�  �^�G"u�F�V� ;F�r�F�( �G�G"t�^�&���^�&�G*�^���G"t�^�&���^�&�G*�% � �F�Ì�;F�r�F� �F�V��F�V�~� u�� �F���F�V�9F�s�^��F��v��F�&����F�-��Fڃ~� t/�v��`�^ԋG
�W�FȉV���^��F��v��F�&���~�r��^܋F�&�G�F�V�F��V� &�G&�W���F�^��v�Ì� RP�v��r��^�G"t�^�&���^�&�G*�^���G"t�^�&���^�&�G*�% �+F� �F��F�F�V�F�V��FЃ~� u���n� �^� �FԉF̃F�3�t�^΋G
�W���N܋^ރ�f;�w(�^�&�G���^΋�F��tP�S�^΋G
�W�F܉Vރ~� t�r�� ^��]� U���V�^�O"�G�W�F��V��^�&�_O��&�  �v���+�P�^�G*�P���v� P���v�N��u+���v���t�^�g"�� ^��]� U����F�  �~ t�v�B�t�^�O"�^�G"t+�P���v�Z��u�F� �'�F���]� �U���WV�^��F��F�^�G�F��u� P�M�^��G
�W�F�V��^�&��u�_�v�&+w�~�J�u�v�Ì� RP����u
�^�&�G�6�|� �^�&�_
�~�&�E&�U9u9Wu��&�_
�F9Gt%�v�^�&�w&�w� P���^�&�G
�u+��� �^�&�w
���^�&�_
�G
�W�^�&�F��V�&�G�F��e�^�&�G*�P����u�F�� �|��^�G"t�^�&���^�&�G*�^���G"t�^�&���^�&�G*�% �Ì� �F��F��^�F�&9Gw�[��^��F�&9Gv�L�u��v�Ì� RP�^�G"u�c��^�&��a��F�3���^���o�^_��]� U���V�F� �F���F�����-<\t6*�P��t�^&� t"�F&��F�^�F&��F�^&��F�
�u�� �^&�? u����v��P����F��u�+�^��]� U���^&�?\u!&�\u&�.u&�\u&�.u� �+�]� U���V�����J&��F��V��F&�w&�7��F��v��v���F���^��F�&��F�^�&�? u�V�| P����v���P����t+��� ^��]�U���
�^�G"t	�^&�G��^&�G�F��v�v
�v��F�t����^
&�G�F�t&�O�F�V �F��V��^��F�&�*�F�=P v-P �+��F��F�  �	��	F��^��F�&�*���	F��^��F�&�*�	F��^
�F�&�G�F�  �^��F�&�*���	F��^��F�&�*���	F��^��F�&�*���	F��^
�F�&�G�^&�G
&�W�^
&�G&�W&�G����]� U��WV�v�~�� t
�� u+���� u��� t�� t� ^_]� U����^�G t+��A�^&�G *�" $��F�&�*�+F��F��F�ÌF��V��~�|��^�&�XAu�&�G% ��]� U���WV�^�G�F��u� P���^��G
�W�F��V��^�&��u��F&9Gs� u!�^�F��� �����ڹ ��F�� �^�&�_
�v�&�D&�T9u9Wu��&�_
�F9Gt%�v�^�&�w&�w� P���^�&�G
�u+�� �^�&�w
�7��^�&�_
�G
�W�^�&�F��V�&�G�F��7�^�&�G*�^���G"t�^�&���^�&�G*�% �Ì� �F��F�F9F�s�^�G"t��^�&���v�v�v��v��,����F�3����^����^_��]� U����F�V�F��V���^�&�*�ÌF��F�N�u�F�+F��]� U���LV�"&�&�W�F��V��^�&�$*�P��F�P�F�P�^�&�w�4��F��u� ��^�G*�+�W�F�V��v�RP�H�F��V��v��v��v���F��^�&� t&�w&�*�% P�(���^�+�P&�w� P�0�FމV��t� �v��v��v�� P�h�F��u�u��؋G
�WF��F��V��^�&�G
&�WF��� ��� �FމV��f� ��F�+�)F�V��^�&��F��F� t&�w*�% P�v��v������v��v޸ P���^�&�G�^�&� t&�G���+�QP� P�w���^�&�G&�W�F�V�F�+�F�V�F�V��v��v� P�d�F�V��v��v��v�� P��F��u���^�&� t7�~� ur�~� s�F��+��^�G
�WRP�^�&�G%? P���+�F�V�^�G
�W�N����F��V�FދV�9V�v�-�r9F�r�#��~� ur�~� s�F��+��^�G
�W;F�t�� ;V�t�� �^�&�? t�� �F���V� �f� ��^�&� t
&�g�&�G@�F���V� �f� ��FދV�9V�v�p�r9F�r�f��v�F��V� �v��v�� P�r�F��u���؋G
�W�3��^�&�G*�P�^��G"t	�^�&�G��^�&�G*�P����t� �^�&� t&�G�^�&�*��+�v�F�Ì�ƉF��^�G
�W��;F�w�.��^�&�? u�"���P�Ì�! RP&�G *�P� P��F��V�@RP��P��F��t�= s�}�= w�E�= u���j��v��v��v��t��t�W��^�&�u�>�.u�>� u�<��>�.u�2�&� t&�G� �^�&�*�+�+F��F�V��^�&�G&�W�v�Ì� RP�v��v��P�����t�6��6��v��v��^�&�*�P�}��^�&�G*�+�&G&W����+�^��]�U���V�"&�&�W�F��V����J&��F�V��F&�&�W�F��V��2&��F����t"�����F�V�����F��V����F���v��v��W�F��v��v���F��6&�? t������^�
G�^�&��F�&�G&� u
+�&�G&�G&�G  �^�&�? u	�� �F�^��v��v��v��p��F��u� �i�^��v�&�G�Ì�@RP��@@P��2&�?uA�F��V� RP�^�G@P� P�2��^�&�G 	&�G+  &�G-  &�G/  +�&�G3&�G1��[�^��]�U�����F��^��"��&�&�W���t� �� �9�F��V� �F��V��^�&�G*�� &�G�� &�G� &�G�� &�G�+���]Ð    "  $   &   (   e   f   g   h  ��d  efg	h����� ��  �U��V.�>�. t���y��"&�7&�w�6&�7&�_�F���U.;t.�<��t����.�D�r W.�|��F�7 ��t= u� ���2��_�"&�G&��P� P�X�^��]� UV�;��*&
'.�&�.��&P��/.��..�&�.^]�PV��6&��s.:t.�<�t����.�D���&�.�D�&��*&�'�^X��
�t93�.��.&�>  tG��<dr*<hw&,d���<��&�G&�=&�=.�6�.����[� WP� �.�L2<�X_t�����t� ���� U������J&��F�V��B&�&�W�F��V��$<u� �,��F��^��"��&�&�W�!��t� �	�^�&�G u͋F��V�  RP�Ì�@RP� P�P�> u�X ��Q �F&��&++���@��^�&�G&�G �t&�O��&�G �*�&	G&�g�&�O�^�&�G �^�&�G�^�&�G+�^�&�G�^�&�G-�^�&�G�^�&�G1&�W3�^�&�G&�W+�&�G&�G�F&�&�W�^�&�G&�W	����&�G&�W&�G�ڃ>  t��&�G7&�_9S�5��  +���]�U���0�"&�&�W�F��V����F��V��^�&�w	&�w��F��F�  �R&�&�W�F�V��^�&9Wws�&9Gs�&�G&�W�F؉V��v�RP���F��v��v��v�����F��V��F�+�F�V�RP� P��F�V��F�F܀��F�~� �r�F� ��F�  �^�&�G&�W+F�V�F�V�� +�;�r
w;�v�Ӌ��F��i�~� ut�~� vm�F����F����FЃ~� t��v֋F�F��V�RP�v��v��v���
�t�~� u�&� P���~� t� P��F�F�)F��F�+�F�V��� �v��v��v�� P�_�F��u�� �؋G+F�F�F�;F�v�F�FЃ~� tx�>b tq�F�  �	�F�+FމF�= v�F� � P���P�^ԋG
�WF�F�RP�v��w����F�F�F��V�RP��P�v��[ދF�FދF�9F�u�� P�=��F�F��V�RP�^ԋG
�WF�RP�v��%ދF�F�)F�F�F���+�F�V��f��~� t���F�� �^�+�&G&W+���]Ð�� ��n�� �p�G*�H�� �U���V��� �F��V��p�F��!�^��v��D$&���T&�G&�W�F�%�F��% �&np;F�w�^��]�U���
��� �F��V��� ��*�P�x�F��u���  �g�v�� P�.��t���  �uG�^��G�F��� *�= t= t= t��F�' �F���F�M ��F�s ���v��v��v��܋�]�U������ �F��V�� ��*�P���F��u��  �� �v��v��v� P� +� �RP�#�� �uՋF��V�F��V��l P�F�	 RP� P�g= ��ىN��r P�F��V�@RP� P�I= ��ىN��u�~� u���  �5�~� t�^�&���^�&�G*�F�= u� ��~�� u�� �+��� ��]��U����F�  ��� �F�V����F��V��� ��*�P����F��u��  �1�>  u��   �&��"�v��v��v��6 �v��v���� �t���]À��  �à� ��*�P�z�� �� ��Ê&t*��u*���� �U���V��� �F��V��p�F���^��F��v��D��&��F�%�% �&np;F�w�^��]�U����� ��*�P���F��u��  �}�� �t= t$�i�^��G"t� �� ��*ɊG#*�ȉ �R� ���F�� *�F��~�u�^��g"��O"�g#�*�~�u�~�u�^��O"�G#��   ��  ���]�U���V�� % �F��F����   ��  �� ��*�P�G߉F��u���  �<�v� P����t���  � �> u�X ��Q �&� �&&�W���������� ����RP�Q��"�&�&�_�������@�F��t
��� ��^�G"$<�A�� �~� u��^��6�&�D�&�D&�T�G�W�v�t��� �G�6�&�D
&�T�G�W	�� P�ƌ� RP� P� ً^��G"u�^��G �^��G"t
��&�G���&�G�^��G�6�&�D�G&�D�G&�D�G&�D �G*�$�@�F�&��Όƃ�!+�*�*F��G:��; P�F����! RP�G:*�P�؋F� P����! RP�^��G*�P�s؋^��G*�F��� �F��~� t�^��?;uD�^��F�� �F�  �~� t8�^��F��N�(G�F��N��t"�
 �f��^��F��*��-0 �F����F��N�릋^��F��G8�G:*��+�; �F��6��6�SP���+�����^��]�U���
V�� ��*�P��܉F��u���  �N��� �F��V��^��v��D$&�GVRS����^�&�u$&�G&�W�F��V��^�&�?	u&�t�ހO"^��]ÐU��~�r�~�v�~�r�~�w� �+�]� U��V�v�< t�<.t�<;t�*�P���t�| u� �+�^]� U���WV�F�N�u� �^
�F
�*��P���t�^
�? u+���F
�*�ֱ����^�F&�*��P�O��t�^&�? u+���F&�*�ױ����� r	�� r�N;�ts����� ��t�h��^
�?�@^_��]� U���v�v�v�v�v���P�6�]� U���V�v�F�V
�F��V��FF�V
;F�vYV����uQ�FF�V
H;F�u;V�u�*�P���t�^��F�&� ��^��F��&�F�D�*�P�k��t��^��F��&�뙋�^��]� U��V�v�v�v�� P� P�Հ<.u�< tN�^�F�&����v�vV� P�=����F�D�*�P���tFV�$��t�<.uF�F�V RPV� P�	�^]� U���V�v�F�  �F�V�F��V��v��D9F�s'�^�&��F�<?u� �+�	F��~�?t�^��F�8t�D9F�uD�~� t6� �4�^��*�P�q��t�F��F��^�&��F�<?t�^�8u��F��F�델 �F���F�  �F�^��]� U����F�P�v����v�v�F�P�:���]� U���V�� �^�G$�D�F
Ft������D�D  �F�D�F
�V�D�T�F�V�D�TSV�OՀ|�u.�D �t'�|u� �� P�^�G��*�P��= t�� �+�^��]� U���v
�v�v��ԉF�V�v
+�PP�vR�v�P�]� U���V�� �^�G$�D�D  �D ��	���SV�Ԁ>�t� �+�^��]� U���V�� �D  �^�G$�D�F�DSV��^��]� U���V�� �^�G$�D�D  �D ��SV�Sԋ^����G�W ^��]� U��VW3��>b tO�G�>�  uF�� �g2�	� u8�~ u����6� �6� �6� �6� �3��拌� ����tQV�6 F��r�� _^��]� RVW3��>b t�H�>�  u�� �g2�	� _^Z�U��VW�v�^���扜� �D�� �g2�	� _^��]���  �K/G0G0G0G0d/j/G0�/G0�/�/�/G0G0�/G0G0G0G0G0�/�/G0G0G0G0�/�/G0�/G0G0�/G0G0G0G0G0G0G0G0G0G0G0�/&0G0�AAAAAAAAAAAA��� ��	 ���"#_#_#_#�#�$�$�$c%o%p%�%�%�%�&)�P�
��*X�P�
��*XÁ>��u��>&�E��������� ��>��/= u&�  &�E  &�E  &�E	  3�������� 3�� 3�� �   ��  �� ��� ���� �� ��@�� ��� �S�� �l�� �� ��>&E&U� À>� t%�>� }3����>3��� P��/X�D�Ë��V&�?t&� u	&� t노 ��2���.���.�U��N]X� σ&�=  t�Ü��u�k���u�	���uT��<w�.�>�. u���.��.��.��.�؎��м�����&��&��� ��2��.��/.��.�&�� �]�.�.L2</w��R��� ��^�.��.�؎��м������&���=��t=  t�'��� �%��� �L��� .��.��&�
�����P�  P���^t�D�Ș� VP�@��ȋ� ��2�.���.�� ���� .��.���&�6���
��� U���~����/��]� .��.�
�� �� �� � �6�>�&�.���U��P�F
��F��F��"&��&�G��
X]���6"��D.��.�� �� �� � �6�>�.��
�     �>b t-��v�> �6����) )p�p�n)G��%���Z�.��.���� 1�!    ��`t.�.�2P.��2P��=\\uY�}.\uR�}.uL�E,@�e��ASQ.��.�ۋp�n:Gu:g$t��%���@Y[
�t��E:\�E �E  �E  �-�X�   .�3�<3P.�3.�3.��.�6�6��6:.�3�SQ.��.�p�n:Gt>��%��Y[.�3��3P.�3.�3.��.�6�6��6�.�3˜U���F]���Y�66� [.�3��3P.�3.�3.��.�6�6��6�.�3�U.��.�.6�F �����F]�.�3�.��.�؎��м����.�3��=&�, �I�!���tP� ��PR��tP� �8��������J�>�>\ t�!5�!�Ȏ�.��2.��2��2�!%�!3�3Ɋt�u�TSQP����VP����:��	P3۹ �>�!C����:�o0PS� ��U��/5�!�v��D�/%�V�!��]� U��F�L�!��]� �=#t=t������.��.�؎��м���>� t����_=  u�^����.��.���&�6���
� �����?�!r����t������IuP���X����rC<u����r:<
u����r1< u����r(< u����r<mu����r<su���r<gu���r<"u����r<"t����
���r<$t<"t���2����U������ =�!rZ���F�  �Z�؎��M�rG�m�rBS� �F���؉?[��r/�F��~���2���~�uӿ�R�~�~ʌ�>�>�!�  s� ��]�&�, 3��
�u��
�u����� ���  ���ôR�!��&� � ��������� �$�(�,�0�4�8�<�@�D�H�L�P�T�Xô0�!��=
r�> wt	���P� �< �
G �!�#�$�&�'�",�&6�*K�.��2m�6r�:t�>��B��F��J��N��R����P� �/[<�u,����t&�3��/�� u�3ɆϡRSQP���� P�E��U���� =�V�!r*�F��� �D�^�� ���!r�>�^��!r	�����3�3ҋ�]� �>\ uø�:��4PS���� /�!S� �_�!� O�!� Z�!�>^ u� C���!�/%.�L2�!�>^ t�NP�c��� P����6F�Q���U���V��� �F�V��&��� ��� &ƀ�  RP�ɋF�V�F��V��	�~� u�F��^�&��F�
�u��^�&�? t�v�����W ��^�&�?/t�x�F��^�&�*�-D = v���.���9�F��^�&�?:u�F��F�  ��~�9w#�
 �f��N�*��-0 �F��F��^�&��F�<0s׋F��d�� �F��^�&�?:u�F��F�V �F��V��F�  �*��^��F�&��F��~�s�^�&�? t�&�? t��F�&����^��F�&� �F�n� �F��^�&�?:u�F��^��F�&�,A�r<vr�r �k�`�#�\��Z��5
�t�6H������b�F��<�^�&�*�P�6J�����9�9�9�9�9�9�9�9y9�8�9�9�9�9�9�9�9�9�9�^�&��F�
�t< t�<	t�~���6L�W���f�+�^��]� U����F% �F��v�v� P��ƉF��F��V���]� U����F�F��F�  +�P�v� P�w�F�V��F��V���]� U����F��F��V�+�P� P�KƉF��V���]�U���V�>\ t��3�� ���2�� ��RP���6�6���w�+ƉF��F�P�>b u,�F����@��6�6�P�����Ã� �j�l�"�  �6�6�)��N�+��ډj�l�j�l% +�jl�6�6���RP���� ��6l�6j�������6�6 ����j�l+�ډ����+�P&�w� P�?ţf�h^��]�U�������j�l+�ډN��^�N�� ��rw�t�62���� P����F��F��F+�jl�j% �F�jl�f�h9lrw9jr�62�>��� P�x��FF�v�F���]� U����6l�6j����F��V��F+�jl�j�l% +�jl�f�h9lrw9jr�64����� P���F��V���]� U����Fz= @v
�x�z  �^�x�G�O�� �z�F��V��Fz�F���]� U���V�n�����F��d9F�v�F��d��F��>b tY�d+���@�� 9� s
�66�)���� ;� v�� �� P���t�68���� P�B��� ���F��F��d�V�f�h+jl�F��V��>l
ws	�n� ��^� �~� |�~� u�62���� P����v��v��P�M�F��F�;dv�d� � �& P���� ���F�V��6 �!�>b t
V� P���� P�-��D
�T��� �&  ;�v*�D�D � �& ;�v��F�V��D
�T�F���+�P���^��]�U���
WV�>b t3�6�6����6�6������+��v��  �� �F��V��#�6�6���j�l+�ڃ��� �N��^��f���v��v�� P�!F��>Z u� ��>�F��N��F�  �6�6�H��f�h+��+N�^�SQ�6:�J
��+�P�6� � @P��RP�6<�0
���6�6>�"
���/��v��v��������+��RP�6@�
���6�6����j�l+��SQ�6B��	���v��v��6D��	���F�^_��]ÐU����p�F��&�^��G$*�P�� P�G*�@ P�6*�	���F�%�% �&np;F�wʋ�]�U���V�F�  ���F�V��F�  ��F�P�6,�O	���^�&�G �F�F��n9F�tP�F�P�F�V� RP�H��F�P���F�V��t��^�&�G*�F��^�F�V�&�&�W�^�&�G�^�&�G롋F�n�u�6.����� P�����F�V��% �&nP����p�F��� �F�  �� �^��v�&�&�T��W��&�W+��F�V�^�&�4&�DF�G�W�v�&�4&�DF�G�W
�G �� P�F�V� RP�h��^�+��G�G�� P�u��^�G�_Ǉ�  �^�F��F�G$�`t����G"�`$<�A�O#�G  S� P����v�����v� P� �RP�I�F�%�^�&�G&�O
�t���F��% �&np;F�v���^��]�U����p�F���^��GGt	�_&�GC  �F�%�% �&np;F�w؋�]�U���V�;�F*���> u�X ��Q ���&&�W�F��V��^�&�GC @u���#�F�
&�8Fr��60����i�� P�I�^��]� U���V�&�&�W�F��V��.�0�F�V��r�F��^�&�GC��+�&�GG&�GE�|&�GI&�_K&�GM  �>  t&�GQ ��&�GR&�_T&�GV  �p�F�� �Q �ȊF�*�؋���F��V��^��G�W�F�V��F��V��^��F�&�\�^��F�&�\�^��F��v��D@&��^��F�&�.�^��F�&�\�^��F��D$A&��^��F�&�.�^�&� �^�&�GO ���w�wR�v�> u�X ��Q P�1��F�%�% �&np;F�v-�F�*�P�X��F�^���v����D&�G�> t���X ��^��]�VW� =�� �!rM�ظD3ɺ� �!P�>�!Xr9
�t5�F�g
�u-<2r)�@�g
�u!�A�g
�u�� �B�g
�u�� t�� 3��� _^�U��VW�C�^�g�� 2�_^��]�  U������F�V��^�&�G&�W�F��V��£��F�-	 �F��V��^��F�&�?�t+��$�^�&�?�u�&�tu�Ì£���  � ��]�U���V���F�V��^�&�G&�W�F��V��6�F�F�F�F��F��V��F�  �F�d ��F�  �N��N�~� t�^��v�&�8��u��F�^� u؃~� t�F��^��F�&�?tt+���^�&�*�Ì�@�N��^���;�u�;�u��F��F��������F�&�?�uŋF���&@@�:�F��^��F�&�?�u��F���&@@���F��V��F��V��^��F�&�?su��^�&�*�@F��F�  �F��N��t�^��F�&�?]u�~� u�S��^��F�&�?Xt�D��^��F�&�?st�5��^�&�*�Ì�@�F��V�@�F��F��^�& ���F��F����^�&�?�t����^�&�?�t���� ^��]�U����>\ tH���F��V��^�&�������F��V��^��F�&���^��3&�&�O�F��^�&�ˋã��]�U��VU�v裹�ȴ@� �V�!]^��]� U���VW��F�  �N�F�V
�~��
�t��
u�y�-��F��ۃ� �ڋ��3��t�����0<9v'��F����u߈O���D�O;�r��F�_^��]�  U���WV�v�~�F�  �F�  �F�  �v����=
uG�F�
���=	u(G��+F�F�@% - �؉F�F��N��u�� F��=%t��E*�=f t#v�Q=% u�D=c u�,=d �^�F� G���F� ���F� ��~� t(�F�^�G��W��F�V��t2VR�v��u��v��v���F�^�G��F��tVP�U��v��)������ �~� t�F�^�G��F��F�^�G��F�~�s�0F�~� s�0F�~� s�0F+�P�v�V� P�D���~� t��:F�F��F��F�  빀}du�
 �� �F��~� t�F�^�w��w�VP���e��~� t�F�^+�P�w���F�^�G��RPV�v��҃F�^�G��F�/��%��=l u���=r u� �=s u���=u u��=x u�o��G�F�F�  �F�  �F�  �= t��� ^_��]� U����F�F���QP�v�FP�����QP�1���]Ð      caBuffer�� � �      Drive %c: = Driver %s unit %d
 Device driver not found: '%s'.
 No valid CDROM device drivers selected
 Not enough drive letters available
 Insufficient memory
 Insufficient far memory
 Not enough expanded memory, reducing number of buffers
 Expanded memory allocation error
 %uld  bytes free memory
 %uld  bytes expanded memory
 %ud  bytes CODE
 %uld  bytes static DATA
 %uld  bytes dynamic DATA
 %uld  bytes used
 Usage: MSCDEX [/E/K/S/V] [/D:<driver> ... ] [/L:<letter>] [/M:<buffers>]
 Expanded memory not present or not-usable
 Illegal option '%c'
 Illegal option
 Cannot share drives
 Incorrect DOS version
 MSCDEX Version %d.%d already started
 MSCDEX Version %d.%d
 Copyright (C) Microsoft Corp. 1986-1993. All rights reserved.
 Unable to load translated messages
 
�  �����������������3�   a    ` RB�� �  ��� ��O���� P�8 PˌÌ�+؎�� � ���G����+�� �������t	��+Ўڃ��������t	��+Ў���N���F��$�<�u����<�uk�¨t��-� �3ҭ�����Î�������t&��� �t�� �܌�@����&H����Ë> �6
 � - �؎��  ��֋��.�/�@� � �ʎں�!��L�!Packed file is corrupt
 %�%�%�%�%� �6�>CC                              ;
;    Translation:  USA
;
; File MSCDEX.MSG -- Message file for MSCDEX.EXE CD-ROM FILE SYSTEM
;
;
;**************************************************************************
;
;  NOTE TO TRANSLATOR: TRANSLATE THE INFORMATION BETWEEN QUOTES " " ONLY.
;  If more than one line is needed, begin the next line with db followed
;  by the text between " " and end each line with 0dh,0ah. Thanks.
;  Do not remove or translate %c %d %s %ud %uld %d.0%d as these mark
;  replaceable parameters for MSCDEX.EXE.
;
;  Use the ';' (semi-colon) character to mark non-message lines.
;
;**************************************************************************
;
;
;
; msg0 db "CDR100: Unknown error",0dh,0ah
  msg0 db "CDR100: Unknown error",0dh,0ah
       db '$'
;
; msg1 db "CDR101: Not ready",0dh,0ah
  msg1 db "CDR101: Not ready",0dh,0ah
       db '$'
;
; msg2 db "CDR102: EMS memory no longer valid",0dh,0ah
  msg2 db "CDR102: EMS memory no longer valid",0dh,0ah
       db '$'
;
; msg3 db "CDR103: CDROM not High Sierra or ISO-9660 format",0dh,0ah
  msg3 db "CDR103: CDROM not High Sierra or ISO-9660 format",0dh,0ah
       db '$'
;
; msg4 db "CDR104: Door open",0dh,0ah
  msg4 db "CDR104: Door open",0dh,0ah
       db '$'
;
; msg5 db "	Drive %c: = Driver %s unit %d",0dh,0ah
  msg5 db "	Drive %c: = Driver %s unit %d",0dh,0ah
       db '$'
;
; msg6 db "Device driver not found: '%s'.",0dh,0ah
  msg6 db "Device driver not found: '%s'.",0dh,0ah
       db '$'
;
; msg7 db "No valid CDROM device drivers selected",0dh,0ah
  msg7 db "No valid CDROM device drivers selected",0dh,0ah
       db '$'
;
; msg8 db "Not enough drive letters available",0dh,0ah
  msg8 db "Not enough drive letters available",0dh,0ah
       db '$'
;
; msg9 db "Insufficient memory",0dh,0ah
  msg9 db "Insufficient memory",0dh,0ah
       db '$'
;
; msg10 db "Insufficient far memory",0dh,0ah
  msg10 db "Insufficient far memory",0dh,0ah
        db '$'
;
; msg11 db "Not enough expanded memory, reducing number of buffers",0dh,0ah
  msg11 db "Not enough expanded memory, reducing number of buffers",0dh,0ah
        db '$'
;
; msg12 db "Expanded memory allocation error",0dh,0ah
  msg12 db "Expanded memory allocation error",0dh,0ah
        db '$'
;
; msg13 db "%uld	bytes free memory",0dh,0ah
  msg13 db "%uld	bytes free memory",0dh,0ah
        db '$'
;
; msg14 db "%uld	bytes expanded memory",0dh,0ah
  msg14 db "%uld	bytes expanded memory",0dh,0ah
        db '$'
;
; msg15 db "%ud	bytes CODE",0dh,0ah
  msg15 db "%ud	bytes CODE",0dh,0ah
        db '$'
;
; msg16 db "%uld	bytes static DATA",0dh,0ah
  msg16 db "%uld	bytes static DATA",0dh,0ah
        db '$'
;
; msg17 db "%uld	bytes dynamic DATA",0dh,0ah
  msg17 db "%uld	bytes dynamic DATA",0dh,0ah
        db '$'
;
; msg18 db "%uld	bytes used",0dh,0ah
  msg18 db "%uld	bytes used",0dh,0ah
        db '$'
;
; msg19 db "usage: MSCDEX [/E/K/S/V] [/D:<driver> ... ] [/L:<letter>] [/M:<buffers>]",0dh,0ah
  msg19 db "usage: MSCDEX [/E/K/S/V] [/D:<driver> ... ] [/L:<letter>] [/M:<buffers>]",0dh,0ah
        db '$'
;
; msg20 db "Expanded memory not present or not-usable",0dh,0ah
  msg20 db "Expanded memory not present or not-usable",0dh,0ah
        db '$'
;
; msg21 db "Illegal option '%c'",0dh,0ah
  msg21 db "Illegal option '%c'",0dh,0ah
        db '$'
;
; msg22 db "Illegal option",0dh,0ah
  msg22 db "Illegal option",0dh,0ah
        db '$'
;
; msg23 db "Cannot share drives",0dh,0ah
  msg23 db "Cannot share drives",0dh,0ah
        db '$'
;
; msg24 db "Incorrect DOS version",0dh,0ah
  msg24 db "Incorrect DOS version",0dh,0ah
        db '$'
;
; msg25 db "MSCDEX Version %d.%d already started",0dh,0ah
  msg25 db "MSCDEX Version %d.%d already started",0dh,0ah
        db '$'
;
; msg26 db "MSCDEX Version %d.%d",0dh,0ah
  msg26 db "MSCDEX Version %d.%d",0dh,0ah
        db '$'
;
; msg27 db "Copyright (C) Microsoft Corp. 1986-1993. All rights reserved.",0dh,0ah
  msg27 db "Copyright (C) Microsoft Corp. 1986-1993. All rights reserved.",0dh,0ah
        db '$'
;
; msg28 db "Unable to load translated messages",0dh,0ah
  msg28 db "Unable to load translated messages",0dh,0ah
        db '$'
;
��2E!����3ҁ*)����i�����& ���� �t�� ��2[@��)���○>�6 P�� -3��� ��֋����.�/�@	�� �ʨ�q�sN�TP�e�c�is L�$ups 0 �y% >   y � !|"U,�,�,�@�<-�-H=� � �� �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         MZ|  ���q/    ��R   !PKLITE Copr. 1990-92 PKWARE Inc. All Rights Reserved    �    ,���@�    �=                  ��D�i/  ; r�	��!� Not enough memory$-  ��-% ���P�#3�W�D��ː���S��9 ڌ͋���������Ƌ���NN��+�+؎Ŏ�� ����u����� 3���� �8�����A����B����H����M����S����g����h����i���r���Jt�s�3�3���Jt�����Jt��Ӏ�s(��Jt��Ӆ�t��Jt��Ӏ�r��Jt��Ӏ�w}.��	��3ۃ�t*��Jt�r#��Jt�����Jt�����Ju����Ӏ�s.��/���V��+��^�u���Ju����Ӏ�r���Ju����Ӏ�r���Ju����Ӂ�� ��뻀���Ju����Ӏ�r��Ju����Ӏ�wE.����t�Z��Ȁ� <�s�M�P�� �����  ����Î��؋ރ���Î�X<�t)�������Ju����Ӏ�r��Ju�����.�����[���3�����Î���&����Ò���ҋ����S�P�Ŏ�3��؋ȋЋ�����      	
                    	
        &���  �	�
��Ʀ�̽�  ����������  �Ω���%   �!$"�#�������'D(  A)�*<+3�,-��.�/0  �12�����45�69�78  �π:�;���=?�>��@  ����B�C��EF��G��  HINJ�KL��M�����  � !#$%&'()+S.�PO356G9:<=>0?ABCD8G41M  NOPQRSTUVWXY[]ab  cdefghiklmnopqrs  tuvwxyz�����  
%3@LZ �d  p����#����͑z�����'5 w ALUc <lu����&� ���0��  �$6CR  [fpy����  ������(  1@KT}��  �� Nz���  ��	4	`	}	�	�	  �	�	
)
K
y
�
�
  0[\ht��  ��������  "'/4  ?BIObmz�  ��������  ��7Vdp{  �����+  :Fhx����  ���-@R �jx������  }#4L]���  ��$7b��  ���!)  059>BFLQ  VZ_ekptz  �������  '6GQ\_io  y�������  ��
&2GS  `kw����� ����%   789:;IJ  ]uv�����  #$;<JKL  YZ|�����  ����� 01JYZ  ~�������   D^}���  $<h����7PcwK  �nx蹘���?�A�: ��9��2��㮉��!   3�RRY�fs��: �+�#���{34��� 4�a-� u�� �U`���&��� ��C��B{��YOS  �Q(�8�0P�3 P�V�6��p@F���S#�`�  A�@���j*t��̡$  ���e���IǬ�S/` ��qd�YX	c*6�< �;\���!��� ��(@OF���"
E�.f5����,|i��D0�-��sN  ��RN���Lřm���?�����  j�u`*�-,Ѽ41�Ğ  c�h����,��%Հ�  ��dY}����A�p��  �?k����hY.��  �Jb�yg��t��  ��EQ�g�
ug�/)G��Z<@6
���0R8g@?H���:�� (ئ̠ݝ� %Aވ�:ZN�0  k�	DjEp�g����G��A��*� �ne|�2���`��� U\ω  ��pe&�̡=�r
  (5L@ҏ# k6�J�Vx���^Y.�>�  
�4-^�vw,�O�  Ƞ���|O�����  Ax�$"���k�l\��4�7gcmd�  *y�0��������  J+d�G�|����� � ]���"��  ����x?��A8�vpuV#��&�
 ��$Ǵ��6 j   �7�-�f�S@�j  ,!�k�!���q�8c � 3!'w��� �Pg�<�dT��
 {��e��"f� <�z�!�N����"�[  �X54p��"���=C'�N�f` -h:��3�nΧ/��
�	;��  ��@��\����1FoW ZZ�7B6���/�!  �E��f�Gu]4  �S8�..�Q�?�p�  Q�<ЇQb��X�FE� ��è�v&LYÀX;J'0)J��J*�k  Y{&l�TpO(-O�LH^  I$�E�<�"�IKѳ� #�6r�u�mzO: ����D'�:H_��  -�^�J�;`��8�  ��))ze�,D@3�NH\ �MI!TA����F�z  7���T��XC�	P  ���y�����IH]� �i1,9�a��% /F�SΡ�7 �C[��p�S�D��ο]& &���b�ތ@�	 �.BI��X��9m]#1����� ��u.c��ؙ1g:�G�!�Qu���c�/J-� �$�〔U-	�8h�<��:�1!p)M/%�
 �i��PdJ��C� 8]Nh�^͒�� p��9��u/� X�0�,_�"� �p�.,^4��:��� �@�Cŏ��9Tp�4!�H0+�', >�L㙍I%{���蠮�<�^ �6E�IP���0L�"j
(� �X���8E�Y�,E������Ix�~Y2�'�A���;�B.x �qb-L�K -_�	A]��=� D���D�H>�^�o0�OAW  ����C��5@�AZ� �9��`�O�EJ	 �W�QTN�!  �F��yG���[�� ����H��  �"p��O2��4g�  �U̣��g`Ǣ���5<�<�� ��eVz*�^+	S �2�e;j� P�j�صAhZ�P�  �C������� ��%N'�BI��;���� 6(0�$���
$  �#��	S���_ �� ��!*p
���8 �
�=A�	#�����)�=`, �]8;��� r�G�C��:�9::�� x�P ma�v�v5@")��.z@��Y�`������H� I-�ש�/�̄^������ )i��*֞ �9*���y�!j.`ŔvfX�W*��dr�YGfe� �C�悝B�.  ��0�����B~d�@@�  +�!�0b�;3,U���z �%���s,��2�" I��"���˘ �1e��<%��B�`�]�j��e; sb�/��hc��V��UY.� V�#��:���: �g�����39X%:�b)�Q  �#� ��tz�U�ee�c  �5܆S�<usJ<0�s�$3k�R���) T�Qᆻ�ȍCu�*�� @�&lY�
�G
#B *�E���"���T�-�	x'��� �i��h28o�N-�2  �=��I4�� ݝ5��0��C�c�^�F���.�C�S��	7���	 Lϡ�`�F��  �5dg�c,W含��F� ���� Xw8� ���1�E<̺[��I �q�y�3.� �����v玙��l �g.�b.f7�^ ¬n�c�
2�] �
3ׯR�&Z�$e$��@
��-2e�Q� ��ۙGC)۞:@S}ŷ2�� ��W�[s(����"/ $]��g�>�p�t(�� [xy�#ʱ Bq�J�qt�����k @��A�S��C}�o*k@�s�'44|�  ����',��h. @V���*����ާ�6 �� �� ��p�P� b��L�/�  @,��c�ChE���Q�h�|�)@�>@<��!  �Ubh�B5#�� `�e�9�����	������T� ( �]��u�<�*�$��" �#����  TE���G�F�'�e�  ��	�h�]0�jdn�� �p���Z�����  ��`�kBc(߬F͸p� 72@W���X�MEl�  �y���'�@8�p #g� ��EP���6u�yV�`� >�/G>� @J����6��O(�(�` �[����ȁnh+U�$��8-�6��c��0&uC@g{kEKu� r���lAD "�M/h�@�Ƥz2@�"( T�BQ��L ȴ�jFE�E5�ߑ �@ �lڊ��%`�  �O������HƋ&0 -��YwDY.���U �:��jC���,� '�dZ`*�U<�#@9P ��[���� *����"��6` mEPY3bw�UȪ8ZGh�&�M��� [��P'�o  ���=`�T�k7k  �Ǭ���"��'�'��  p	fi�j� 0ǧ8[� `.X[}ѐ��ata  ���~��)d��  �r��C���3  �N�����������~D�� <nk�j� 瑄6���� �%UB�3��K"� �뗯0� �Q�n� 'p��;~�< e�G��X �Y.��e�� p5k�lG��`�Dj��N�[X  �Vڈ��5���:  �o�h&�F q����d0 w��4&�_�}!d� ��b��d�#}�9��
>��� U	榲��=}�  ?Dm��i��#k%�S@̰d��� �?�v�v���m�<�����L�  ����
�*Dᡎ	g ��X��\��@�(�̱U�1"g z�RR$:��\?g��t*��������x -��`�?�+��� V�Yj����n�j  �C����P���, F�����9��F���#��," �����  Hi"Г`"��( ��(��C�X�w  J�:yZ���8^JW ��$�EN�lN�  ��P��H·LgM��� ��I$P�=�y�t[XJ@�����\CJ쯠� ��|�7�8�o��`�T��O;�\��� ��IS�	�	/e#  ��ۨm��P�$��2�  wާ�	�5��Ax.  �z�)�f 	���;y2��T� @gX	-�� �Uc� � ��͜�t
&�(�,���C��:"A d�� ��9Z�u~Y�h?7n��$�k�����_� p/�'�(�� -
 R"�G'�, �����ʁ�� �8Y8wt�p��H2��- Bzt$�°j�O*��+r(` (��$�n�����"  {��#28a�������� � b' �7|�+	>�� �DsB!D��3 CW�BS��� �Qٙc $Q*�DA4 B!q��J��a# 0�x �����  /Yb"
�N� :�,��A9� ))Y�W�����D� "��Ib$�;�E���{4>Hdp�"LEX���S�@  ����Q+��h!e  8�� �q�qyN�@�������	�&��jI�d= -O�%`�1P�" Y������(1������Dp41�#  s�A���  �)���?H�h{P�X��$�$�<��S�$ay�� ?��@D�f�ӶN  i'S���?���p
�-"� s���P8�N^��� 0#hv�S��:*�r n��� �<�@ �B65VS�uIEu  ���8�T�����uIHI�r=ࣰ��}�q|	�%� @�����'l��N�"�1O $��by\ )à]�1�;N2�����+eI�]jy�*8>%���`@�d��b�e�2
��}�pGQ �����I����V:)]�)YE].\ ��1�5�U  �3�+�#K/� �"�����;�f�m= ���'  WF�_��Q�K�  ��,ݑ�,C��n�  (�.,zu����(�Ai�  �	���CLo21E�m7�#/,��� �v��4i�Bj�Qx@f�{�� D*� hp֛���pE��5 ����@<b�d�v  ����wx�XwhK�aPQx�Q�4� :�W#I�x�נB"��`���x�Q=&�h?��i1�����e�dO��4���>��b޹��
�F�^#Td9�g2KJ(��y���  alt�G�����* ��,;�,�YN8c� ?- �(�ûC@
	���
{������)^�S�!  -�=�qCc��))\)�~���%�h�8t" ��Z��ĵ�G�# 4p�/f˩�kZ  *� U��F� ]�   VW�N�����   �u
�6�6�HrM�� �
 �� _^��;���~�v ���P�F��M�N�|  2�  �³��B�����  혓^�/tF*��� x�s	�늇� ���+0���XS��][ � �QB.EXE LIB=�lQLB d&�<y� ��� NULL STACKYMBOBC_SA0	 � B_VARSN �  ��y��Y ��a�_�\�] �X�W P�R �.9 �S% X` �! �>�{t���.�>P�u*�;X�"�L�!����  �����qt ��2����� ��	��д4�� �������:/\.�ǁ�0 ,t*����3�QW� �O������uGG  �;�r�_Y��w��;�  t3�[8Nu�f�� ���3+ȃ�v� ��l��u���c��I���Â����6˴����7аJ`�� =�ô>� o�����V�v  &�
�t#<\t</t< :u��V���1 r �R�����X�d�c �V�APA��D :\��ZB�G[r` 3��vPS�I (�u0���7

��t3�`$SRP� ^]�  @GI�~
���I�N���W����v���3ɶ
<;  t�A����3��AN�谌\:����:0t�V3
;� ������^s�ҁ ~Gu���9Fu�� C�������_��
 �s6�} &,3�3�II�t����&8u�& R�==u�G��<' l��(� x�(��(��(d
�ǌ
�(t
�(��l�)�!�` U�ٻ2� K.�!`�.�&�.����]r� �b��� � ?\=��
 t = vP�ZX-��u0�������u�ħ��
������ l�@O������6@ B��PLOO �RPDF Tr � 6
 ���BBJf�� *���RB��R_�_@PE��B@@9@�@�BPnO Od8r��4�T�y(B8?K5?OS�3h Ԭ �d2 ��4 �S�) 	"9"�/	Xb��� ��{W3�  �N���~���s }�_]�@������ަ�~�%.�,����;�s��	�0<�ح;�A�;�5u�����^�V `��߬�'C#�:����@�rtHHWQ ���X+��&�_��Wai��+��*_  �[XSP�Uc�R�Ý�^�*�����	+s|�+�N�E�H������@�^M�S�V�@�! ��s�9 �l�`�%�o��(��隴<it�����o j.;�1 X"�Ѐ3g�
=��= u��[� ��0  ��q(�r�3ɇ~6�-�>�-'-lc���ѴvF/���6���P�b�p��6��-��n�a�R�v��1([� �[# �G���uF�6  �(�tNNV��s�� �@t�L-&�\S��T��.�H�'�,s� �ˋ�=3� �h ��� �tS�^! ��t a�.f��-X�>�-��-����X�&�-��PQ�� IIQ���YX�=�(�(�4�s��+
�"�E5.
;�����Y��
Q� v�� �������-��Q���Y��
�?�V���؎��Dڊ�2��������A������ &�~,� ���،��󤬨t�$� �^�{+&���t�@�*�����Ȁ ��&���2�Y�� S��PS�4r P�q� ���[  6r�[���7[X��� `����t�7�_�04+��X<�i y0��h ���'� t<t<t0�n  1���5�1Rj�ii /: r�G��X@��&�@�mJj5�  d5��R7+��a-u��e� �F|�8	VW6���%3 ����]F��l\�8^��9Zu���&&�q��96�u�]N< N�<H���.��� %7�  �uրN�����u��~������ÀE�a<��&��4�� �4�4먃>f5��=�s뛋��&<�� ���� ��v��+��P)��� f�
 �>���FF%�V  �u�H6�=�(B�>6r@��0��@�]�- @$A���X6y�V%�M�������V��6>��
��� P@�#�Q�+��3�Y��X����h�w�P�
�f�F��RV��R)D��v�3�6 �b-�3V�34�'�s t�?u#-KK�r@��G��q�3��3+�]9-t�7�?u=�6���7?��u	�a3W�"�N3�%P�d��� ��Q�J�����$��@�@�9�X�5��W�03�*�v�..�����FHFHtAA�� �����R���2��2pA: 9��a	 0�} @VGK�II<t$< �t���.������< S�K�2X�/u���R�� ��1`�C=�ЫwJ&����G�����u�΀1�uTR�d�j�Za`@�ʡ�R��]���K2�H��p�V���r�E2��ZPP�����2��+�P;$H�t� �2�� :���I�8 zz@�2`��pq�?{�G�O ���x
�LtJN +�m+���� ��
=��v�a�
tu�  
Gu#�G�ӡr@(G�r�(w���K���3� ���3�����r ���1���r(�= Gl���u�Vt����c �� �k ����"U ` )�N���rF��0 3t�� |<�a&=�U!18�/n�l�, ~'��<�dw�<Q�H��E���3:I �������r4t
�1�@����(�r�\t%Iu�< ��L ����0�F�0�0� uF��sBU��$�$�3.�3g�C4�1�@θ` N!�X�^mK����P+���P��Z~	�a�F�M0c��| `�t���2- �|Tx �!�@t,	<��w@�u����;��1@��N�Y_ �68�<vFF����[/��:�l�6\T.l�]ǃ��F� i����<u`T�z����b- �_�� �4H 0&<u��������'<ux�T ���r��]H�� |�~ �t*�����1��@�2� ���keeH��[u[�u�%� �R�`�n�/� �^�����t�`�,*������	:�39<r  �.����<�D����v�d��x�{����u�� '������c�\q�
]W��f�W ��@ t]�>T�'���0�N����4�D���w
.��k+�,%{ ��Q�X� -���N~�t�Ǝ���^|�1��w>J{ �>v=u' hGEue�u��]��t8�� =
 w�� ���d��0p�J!�� ㋇:l�-���-Ou�`��m$�-�E@P�Y>P��-�.y�z�s��	����|�p`u��D -�*ø ��/+M)�''
�{9O��& ù ��!�u�-��3��.�P� 	�]q@u!�`A qt�G�3$s�dq�W9�Z ����4t׸� �V[�F/��0�D�=�%p cDPFE��	D�#	X�~Ԁ#�~�tk6`1.�F�eq=1t����]�u�q�H��f�����U��$�R� ^:��5�` ��A  �E%6��K ��F�T��w
���8
�.� �a)�,'� �	=u�*�t�����B,W�/#o+���	$tk����  |�`�C
�|h�w����Q;&\]�C@�Y��y���.)�+*��u%���}�+V��+-��q��=�EV���-�롷(��� S��+��+ua�F0  ��H�A�k���P(P�+�P�RM ��p-������8��t���*.�6u�w��Há�q �pq�N��-�>b-<s�0�WD�'����%S+�\���u�6����;�1�u6�����l�+�D�� ~�>PZP`����r#�5�2p/�q�o��~zW��* z���ZB
��~�|_�W3�6 ZfUEu$���| c�@��G���� ���It�tRr8C��=À>` -t������ F˰r�3'e,0��X\�*@q<#  	�I'�V�aW�F���-�� �x+�G�F��z�M7��x u	�	AW�}7�A5�,G��5G�|߉��H�>�� �� 
�����ua�?Ұ��DuJ��T�%
�8+pF������p*u/� %(�r���` 9�-t�$qt�W8:P��>f�8�j��+���e��u`<uZCq���uL&r T����u�wz���X�� �'L��C |1t7����;�3y0T! �W��|�+��fq�)0&c�)��L� �`����N1� "�B�~�.4r_K>(K��0��g���`E ��
0	��� Hx�V�\�*��'�q��3������� &	��n#��O�^��&�N� +Ҋ$(�a��V�	�,O
���}��4�*�j�@t�F�
�쳀N��w��* t
+�c��|= ���;Tt.`0,��r!�R���`�dq���8lOr�� u�e+���� 
�  |1�xt��
�>4��X��z|tUF�<1��d
u
��	@��/�}(�`Z��W`3@�{)��: @y6r�� -8��<��s!�	띷�X���5F
r?�����Rb����V4���� Z$��A��? Sk���E	�00%�0��*�~��`>R�$�k�&�����X	s�	u"����|}i���0&�&�}�/�Y��	���6���ր���N�t|� `;�&�t��w�	7� �N� g�|M���n��u�@�	3�r`҉�� BB�rR���|Mz�I��
-��o(� :Ë6�1�"`�)3�\of���(p��DrTX�~e3���s)���$ O�%���8w�UR��Ӏ/�k�t�F�%�Ft۸8�A<%���5��r/�%9�$�a�8
����B|�m%�	�|�Q�1 @ð�
X��ȏ}�|虰#-�����s��_� �` #� @�}ܸ +�����_�<�̐�U
�
�+�`G�]�\q  cq�Xu8��pu�>�c0�
=Mw��6����  =ힳtl �+��  ��� ��&�� �g;�;B�#��&q t�N��g֣V� w	�Ѐʀv-�~�� H�G
*�S�.�؊�r[��[J���!)r�eXeq@QP�6^��Pv�����
Hc'�ko8��+�������t'�f��0�u���?�-T�j& �k��j��4��-�Y-p��Jl�:N��N%�*7{ �<r�n��2r!+�2 �Uu� ���H�c\�)R+�0 D#&�� �G ��@u�^����w�� �� �P�fR̈dD�0 H�t$�� uu�RI���|r�#�7����V���|[t
_0Z ߳�:��*u*��o�[�2J	 ]	 ��eq �6bq܊����"���"��"#�Ѱ�aF�=�V��Pe"u19�MwIr�"��s�"�*�|�?�&Nt
 s�^ø�
D%��i������,D��eG��)	�#᎙�
8r'�Y�Tp�����  Z��|��*,�("�����\Yd ��.ud`���&����d����{ |#tdu/ņ dY�$N��4��63��$+'&��5��E���#P� YtF ]�W�� @;\��t��㽸�Q�FS$��� ��݁�u y 
	���/v������	 v��N,A�< �w{���.��~,������	��.C��Y��Ȋ��$�����*���:�u� nG�r�u1�*�`\�:fu��
ǰ �E��?�t." &�]�u
��#�SY�$�)4V3�� �6r��+f�r/4*�{��x.���b.�<s����i,PE	�h�E4%��(
h������}��& ��"u&�֬<"�t$u�NJe�H3+@ �@� OH���<@
0r.<9w*���P� X"�����rw�0d�*�Uid
_u�N� �r+w���k`�6�����0._�LLP�H�<��\����W�~  ָPR��IN��T��F�F���� �)& +���F���(���$��8��I�G��� !$�r�u�u�'FNtܲ�J�V͸E��V�  <uT��GOuN�~� uH0 �vҬ<���[S�� \�Kt��/�)#�H�0 _�߸�.�Y��N�0 @�V��Asu�g�[�Tn�_�6jϤ��;$<.t����S� D$u@P�m�s	 �tN�p�F�,A�
� ד�N��	��sy�@# ��,<rN�@7I;bE�*E\�-��>
V�@�L���(�̀�^8y)6#��NLC��f�<����.�:	E�޳���M�u��* y�+�l��. ����Nq��
 7�pq��q�� �=Rs���r ��9H-u� �� ���_Ã>B�Gr �v�4=4�@�Ge7�Ǆ�;G���G��3���2��2
9L��x���ϟ�s9N���q\� V�9�(S�K gd�<�H�O�B�X �o+���v�eǥ `+ �5 �����;�W�h�4����v�! �����BJO�%��w��6 b<Q@����%�u�X���@�w�Y�*Kk� ��c�r>t�+
C�r��4�@����@���u
#kw�$�匚uV|���������#SQÃ������>�Br�$ ����8Y��'�X(��s-�g�CQh 3|T�4|O�ny�~������m��-$	� eta�#@���R!6s@p��	�Y� NK��������WR��B�;rwNe�RYxl�\��o�s)}�W� �:��rò�+�PQ)� \p��?���� ��zS�U��"����c�
�3{����<��P��� D�rH-��1Ae8�9��� �K]�y8	���;z_O6���f��S�PRS'\�Z9Xt`׋nl�G���{���V�6�8�;�s��ȭ�ȶ}���b������p(
�KX�G�

AI;�$ +AP@@�.�)f �"  �#��N�J.��� �;&zvߖ�Nq�F ��.�<w1t�a���'?� ��'B:06g�������1�<�r��- ��qG�`<�t��M� �#��ƀ�pv-�R��%�(' =G3- = ��s��-�,����_��-=17���  �|:�X����S�-�U1������|�l�/�>��2�7W�8԰@�\���/"�Iu�6S�$��&!q�\��3��9��&�~�ÐK��܌Z��>� '�0����"]�"b"��� �V>��LEto� r岳��La�t���v ����D���<�0k&�{�؊�#̋����]�����)�#t݋��n�	:�v�߾�!�: ��w:�r		TD��������?|�n��4n�
}�� ����P�4�^�S���	#���r���ƋV�F
! m�s�F��^]N6�<��3�7��Wd�tr�z�q��v#�X��q�ts����f�#��9�9��1z�L'�L�*8���H�� �S�1[pP���^*��j2�f��F���Fn6=��F��F�F�D�|v�!q���*ҁ��+�~� �~�  �<$t%< t�f���  �<"u����<:u�
�u���8��餀N�� Ox���۹���{�C�ܭ����u�~�� H	�n~�����e��gN+�KW�}�N��
m�QP��N����'s@@� �r6rBЉV��]u�S�RĈ܇��H2:u^�� N�^��r0�����v�C����@[��P� O %&!#$"\
	^ �_'()*+,-/:;<=>?��0 �		
� #B �S@oQCCESS ALIA �"ND�!NY �PE1  #SC@v#TN@}�" 1&E 3EnEP�QINA R,GLOAD	 �� ��CSAVEOYVR0�"( 7L	 7o(S	%9πBG8DBL@�1�?EC.CHAQGDIRNzHRD�63T@�W#�E	U ��rEy	0�� ��CLNG@��ۅR	��9��g�%O�%�OM� cMA���D�S
ON!��lST!�!S@�y�lSL�SRLfv@��VD@?S��MBF@�I@�����1�"S� D`�TA 5EE�� g0ҤE)� ��c/EF
,#�E �Ǌ� �F�!?�	�!	�O�!	�!
 	TR! #IM!#�O=QOU7 �RAWY Q{ Jp,�`IF!`,�yC3�cN�R���
D�O v��"QV�GG` 6�� CRDEV��@�D�'R<~��R@� ;R�3XIT�dXP0@ a4IELo�sI�T�@	cGS	� �1�X@p;
I�E@s�"@�wUNCTI�),�8�X  i&T
1#>��d0COS�w3OT�3}lSEXD"{m ߃"MP��K��EYD)hN�-� �UT	�]� �T4�"�LPC�$$T�@FaEGERe ňL�DM�8� yll3Y�|��|0<{ WBO�DPZP(`CC;D]3<�TDd}EN@kT  ?INE
A#�� ;4�� 1I~��eC@tA�W	`��� 7K	cJ�8 $F@{3G@�1�ONG �OP3P���SPR��.�7}������IMD� � -IE���2�����NKDD�]@ Q�SK�D3?�_K(��	�SD�XK��D�"OD� �ơME�wEX�n�T� �P �lD�!FF N	�uN37)	/� � 0�!�R�#U9�0�Q�&���A��c����CC�YN��NK@�%  HA���LAYJ��T#��x3MAP@�GOG`P�?3OKH��WR�E��1��m7
�� /UD)]L7 �)�QO��M �IZQk��ADuCED�Dx�!EC]�gTOj	�6�j WUM�xlTURN	�' oGHTD�C8M{�'bR8���P ����f�'U7Ӭs b �yDD@��]C*NY ��G��� 5 �(A	�G��@LE@�O�M@	�S#GN@	SHv`�D!�IH"LI!		l�v�/�NAL#S��(	Μ�D �!R�C���PA �/	!PC #QR@6OT �ATIC!&1T*�GK@=	3T��l8L��	��?�GAK	?Q
J1�SDR	��B)M�v�WA1_l SY�n � !f�ABdA�Y	1�N��I�E`	rE 	RAd	|O�@POFF�3�ӅYPE!�>�&
�W1�h�EVJT�WNLR�Jl&� d�LS�� �tL@o+AN�RP�v�a	D�	@G@�̜�IES�e���IT	��w��!�CH���IDTH�9UDO.6� !+V � "` OR� �l%Q%�%k  &�&_'�'�'�':(=(M  (�(9)O)�)*"*�*�  +�+,=,s,{,�	�	�  	�	�
�	


%
6  
:
�
�
�
�
�
�
�  
�
�
�
�
�
�
�
 `BT|���!�  !jY"\"V"_"b"" #":���   
����  je����	v  	qNl\	 #x �#�#}#,9?: �2 � �x�  ��iwo�{��n6�!�	(��� � � �=��� � � �` 1�	�# D	_ :Tc`�:���11�	��5�'C^ ��M1<F='	r� �l���
~+KN
��+I%s%�< G' ��9x� e@�. ��#"8�#t8�# (5�(i	nƖ���K�p
B�n� y<m�#����5�� )*+�m,-�>�by}Ry3\3\�d���[�F�G��ԈlH��R^	��PMdJ�R�BI	 Ú(�"��6��Vl�EN,�9Q�&
RP5�O�&0b�9%5�9��<���K�	�TT*/SUz�t�r���1��1�
�;,�SÈDV�ע)aW	0	>��3�C4 �Wc@/��6)��En��h�d"��7���Y�&[�`E�"gGS��g({�	yV� b�&�b�����"�p����i)H� �C e� ���� % ����	PN��O�I�	��4��6XM���V	XG�G��cIsd�[*Tb2c��	d�v��<bY.��_Yj�`@*���r���;e �@=fk�~��)�,��K�W�F�`$F�	Hg��vD"Hl��(� ��3q��།#wD/
��Pm�`�%�g	A
�	дL
�	rxxE.�-\ѕ#<� u��`I�γ��ϕ�k
B�w��\
����/�f'�.�-�)�.��H2L  �>��ޔQ��q����� ͵ co���_�!�hrL/exvl4/w1C�
�4G���E	�%pc4�4*���F�)HFF��(��&<*���J15 L4����(#}#t��Z�:r2o2��G�w0�!��$�{8�6/$3gcu�������19�9b!CM%!6�R(��w
�� ���V2.�	�: ���-z�� ,�3�� D��L��M	j�3v�%��-�"�y"jz	V�1r��1��	��T�$���z�D�O^�3����V{��� �0z�cgo����@cj.'U�	M�	7
4�\.��]�d˽�^N$��{ �� �!_G�������& ��`���*r[,>-Q.m	./��01�r+4�\567.�89��:;r�<=y>���A>�B�ET.�6�F��6IJ�rKL�\MNO.�PQ��RdS^T7UV.�YZ��w[\�MB ]�'��=��]�K�r5��0d� �4p	?�48��� &@F<S;�3s<-s4'h5�	r	D	�DŁQ��� �{ �n�� �@�7� �0�&�;�H�R�Y �P�3,��1�0/KU�)�`�^��<F& *�+ �$�cG@*1Rސv�x�=		2
4Vq	��� M�� cG	]S����r A`�Xm
d �A�.��N'@t�Acg|�D�?�����r������\��e9��!� E��EAg��J��6Ψ7g��  lw�TR\q�b-�F�V�P������ ��v���� .��O��'�� � ��Dt�� ���c��tL�2  �~� *�� �=H r�\
=L w�k�@[��Q2�=Rڋw
��Q@		�d����%aHt��.�����cQ�f
�e��� �=�0�q7���.��~ˀ!�V��t��ҹC�|�~�=����P6������$V+����~@F7 �3�u%�wF� n��X+G<�|�� ��n3Mtb܎͸��t��Z�u��t�� �����Qu��A�N+�N�Mt��;�6� �PQ�Wō
�pfn��c �n��E&CC;8rw���:r�n�NPS�P`��[Xu���2w:��O 1@�V�W�G�����m���t���Xv}��%~>K_^/��v��6{��F�@�� �N�N�A�����G�~ �d�vl���>�:1�(t_ �<tL���1 �l�~�n���<K�Du��f �60>6:`)���0�@$�G�l�%� X���$x �	�������#�+;����tށK��� ��Ei���M�8�q�P<�+��n�F�L�G�X� ���l  ����SP�	]�/��  *^;�s �.���$0 ���7�A.�~,@@�p�.�<���Ҁ~�Zw8���!�� �;�t���֋јB�k�,��.� ����t�$�B��齒�  :� +ۋЁ����u0��r]�&����3 �t�_�Dr(!��j�` ���u
�@u� ��=� 빸�&bz�"�CD�0u u)P�<� �� ����� >�������XPiP�?<��p��Ȱ���� 1 ?��X�V������w��x���V�[3���<SN�):^9�&� ��X�|�Vz�D��O��w *T�Q� ��v��@��u�F��Gx���=�RN� ��6�����<pv�����Tu��보��ǳ������L-��=��T����^r�@6�p  �| ��p���9F  u�
��V�E��+���~��E�|��"� tR�+P���P�;T22��G�D"��CA��aE
D�^�9D �� 	Z8P
c�=�p��8��W �ڄ9Ur���������u�O6�+��ˋN
�>�v�U�3��.��N��64
�y/��Ȃ��`�8Pbq\q  �dq8�0D����gx:��v�����<g�t 0��N�7��E�C@=���+t� �No��� �!Q?yc�>V3���qm�����D�sb�DP�8"u�f��^$OLGr(�E =���s=�	���̍ǵ�u.�G=�L�U�Ac4�^ ����@���?p4+��6�}��>J�9�yu�EӋ�nl�u	�j�fq�+�3�;����G w��v`�[�߆��_[���a�F�B�S,��̃�  ;� w� �#XX ��,��"��
>O�;u���K붳�5�<���u �W$�&�؋v
��&�NӘ&�u��$�#�6 0�-QR�6�->� �t"}f�I�X�P �&��ы�u(QB�D2^�J�W���y `�����;�t#�sxa$�� w�A���p����K'���_��+�+�+����_"G�VP3 m=Rv���1� �>�-�u(X�*u����696�ps��+w��x�S� OO\q���qa��t�3#��5WbqW���� u� a)~��rt �F`�u��\�a8c��2J��$�W�#� t
�t*���N���{���yt7�eq*<��� �<v߀>�o;�u�"? t��xv��΁����b�fqD6���%+�FX����7�	�	t!�]�f��u���'�Y�@͋%�vl�",�MI �u����+]�J�$`q��L���P�	 �� �t4���R�y#�"��ut/a��Z�	%^<��S�$���0�wuF��CC��T�6���p6�"đ@�3$q-$0�����D&q�u�{��9��F���-�~�th�Ɗ��S��
��0��-)3��9s��v��m�-�lN�JT���������t�q�^�0Ħ�G��	F��r�	�N	G�	������#����=��-���,���@��H>�G=�W% �"'bbq��J����v���Gnt
��%O tfv1�x��Ί�,;�����Q$$�>x�D�w�-�J	4fs"E[B0WV�\�>��� :(q���Fn�&���I�bu�De���#�0�F�;u퉥�=+���0�L�@���^_�y��;�z����{��bz��+ƶt�&9-�3q�%�uq�1��v�h�m�D�t��%�s.�;�t� uk$�o��	�L �c��&��L���"�d��]o u8m8''��+9 ��6D����;�t��9D�u�xNyu�h�8�w�������� +xU)Vt0���V� ���f߀~�y��F��؊��iMa�T�W��PO�_�  ��F�^3F�P3�M&��$���B��&�m]r����-r�����g{�?y�������!�^J���z��b���0�j�~�8-�&8�t��-(�yG��yG�;bBԷ� rN���'�a]�]q�2�jC)��t�p���*�� �tT�@A�R,��ta�a]�8(��*23�=�V$I"I�(m�, 5�,�,1� �\6�&e� ��t@��P�c��ƀ�^Ѐ�A��K&<����j3��KN�/DIX� x š�a˚H��u<�t5|�#� v��6� @`��9O��� 2��"�yX �Akusr��K�B>B;k/%�ː�ES��<�@E�G� ~~����^��;pH� tj�d� }uzu�N�"��4
�	Ă�^%�1�� ����(r�l���-�S�
��s�v���r�#�֝�`4�|�	4*ۦ��� �`{��#�Q+",;\
����@"P���� 4G��L$�<���S<��M��-  �.��F�RP�Th�g��� q����O��� $�G��:���T��Eu(èR�����U��w1!)�)u�`N,��޹�E��S�P��U7w4)f���U
3)Q�P�W��#CBT# _ �w
� ��7B��M�F�U�g`�7 -��Mp���e����.�t��e]o�]��G@�L��S��Rtq���R�ه0���
��:�$�P�T�d�t���6�v��"p�3@����(^WN�Ч)G��ܿ���W �����>I�,à
����oq����v�d�~k��E� u�����	uM� tFt ��E�t9�}�t3�E$����'�%|F6E6E����*f�MW'�+H �u���{ݻr}~o����u�@g�F��r��**�$�aj�334�33]���p�uS�$ P��$��� �_t��M�QP�)���V)�73������s"3/�^��-V,1^���  23g�	q�"��	�c���3=\�����G�%�0��Ë&c0�-�AA;<�tًx�V������_�J�Wo����(�L
AttI�u�D�k�Z�h(�;�- ��V���p+�V�S��T����3 �n�ub��t]�t�!�KtRt8�g��G�M%# �6�:��pu x�PQRQ��f � YXS%�0 �2[ �3Z����^�0,r��;n� S�>4:����	�"O.�[����ś������pG3�^"+R�Y&��$�pV#5�"W��)������/��9M�t�e�}�rp���7��1  ����uB��\q�M����@�]�T��]A;�u���"Ph��;�qXt�� �l�ŠC(
1>�{<;��t[S���ȁ ��C�Pu
8���u@u53�w����&<���`{pt#�=u��¶^�%t���=�\���Ru���PFt1'j:��$���| ��BmN8�B�r��\��#�;Tu�
u�S��u3gn7ta�"�� F��ru�l@n��3ҋ�, �,@t��+֋ދO�  w��G�&eq:�t
W��1|
K�������l� 8 8n��@Q� m ��+�PQ��S:�rYfP�O u
�I�l�ދ�BtJl��0��� #�un9�d�(R
2=tc˸��'	��N$��S�ϻ�������~
ij��̃��!��3�o��H��f�M�>b��s b��t������W���-+*HP�|�U��t p;E�u��%'�q;Dd ���������_���Ƌ4-�^�p�+͓�3�S00�(xN��G
Y `HVPW���X[��[V��
���|�oM"�z�� ���L L�����f�@�^���-�>�  ��;�sdW3���ރÈ�L_3���p �D8�"t,	�|���;Btɍ��W����`��
�0W���F
��zu�v�206+0�c�c���	�Ԝ�֣� L����;rIp�H[�� �u���p���
�;	�����=oa����LqP�LP<ɸ@� �gUH�^���PS�T� ���:�D��� *E���~��c��''� /�,#�wO��3*����\
�DW`|T�(r5%�E�?o>F#(�\r�� �<�^oW�S@� �� 3��D�+*k:e{+�.G"�ܚІ�g=������ t�	�h&5Sx �HM��W
�GY��	PR��5ZXˡn���;�t �$�����G
;��u��J���E��"�,>�p�� ��n��� ���p n�pv�&���&\��G魘MAn��W���[�h�@ ��Ǡ�Z[/�R "�  ��߲V2�� Lv�
�y������p�N��Sn�̎2[�I��2�Ci��cK3#���*~����-����D8Mu�� ���&�% G#�:�u���~�ɝ����7"� ?t��T.�`�3��F�J>R &���o�&��t0�f
[4�K��Kj�!��6"'6�-q��#�~f�OȄ����))��� p
���+��t.���_�I�x��&��=}���&�ԋT^׊W�^�sfW�iP�a`�YP����Q�=����&����p���@u+�y�V �)[�G_z\�VW)���_ ~+ɊL����-�X۶�&�\& Q\�X�Q�\Yw��y9v�h&}��@2:�@�	A$�2�<FuO���v	��1��NuG!�����Y�E;�`ɵ�=� �Q2R����3$W��:�[�C
2�
�u�[w)V=�0���� NV��?��䑺Vb�3�5�@��DRu
v� �\^���T! BBx���P�	w��4`��Y�A��f��X+����CN����x�x�)�.�VYU) �����֙@p�� ���>( Y��2��  )�� �Pj�UP��[���;=���X�Q���E��8�!�ڳZ�s3Vq��XDv5VP�|u�zs���i�$�Di��X��%P  ���+ҊT+��B~c�� 	��Z^�� �h��Tw>�-� �-�u�-;6�,6�p��p���z��~y �䞋tFtN�Es�1V��;���v
<����,��t�� ;v�sV� =��t�v�s�m�^s�-�� Z��QN�+�E�@C<���&�p������V ��v� �����_6�����"�f"�`$�^{�Hw| u��m������>�v
�, $G=�F�'[
&dA
���l���Y" n�^˚J X"��-P��= w�P��ӫK }�=��V�����[�~���y"[�pB����Q�����-���,�_�_��{�pt��B<���!��P"=�[��^�<Ww�Y�VE[�4�a,�������k�`0qP
�t0' t2�"��X�"q����9���0x�u��8P��<7�\ˡ�p3 }t	~�p - �~��p��p���!q�A�˃7�P�ڻ 7��#���q
ϡ�AuB��Ɛ,�<��A�A�l ���� �ˋ�� ;�r �t;�r����rV_W@�����2;X�l��?��U���<��P�rt��u�����V�8	v��+����_ջ� S�a.�P��Q��Pٔ����һ ^� �_CtK�G~<M��+*�W�F\r� ��~?F�<(	�h0���  u�V��^�FtE�pNZD؏.;�u�<�r'0�;Tu
�d�[�]:�t�~���)�t����'��.��K��3_A�N�=�P �wX
 xa�PV�
X^{ ��> �\ �,1�EG�����ƅ`�n#����͚��"^_Ë��= 0+�W�����RP8�SQ�� /�E5XXǶwˍ/��\�
*WH������q 4�j�-�G���}�� ��������õ$1�#�J1V�	!1�c	;�p�ࢄ;V;�-u�]��>�g�wn�X
 ��ȇ�O  �W;�t������Twu$1�Su��`�[Za�XqRAO3q�8�j&(ˋ�JBt3J;�uA��N��'"  ��ݾc	h��VW�3�� �~tt	������{κy=B  V;�tC��vb�Fu  \�	�W�	���
 �o���> V��e��&��
�����U��Ep
O'K�$���WD�;�-t(�&�F��
P(����Ff�)���bа �6$�x5�+�'� f�\S�� �ɘP��S��p�&�p���"�qP�G9�$�.�=��t��e��8R�t~��Y�w��u����[P�C�`NG��pc�!�hHt9�FzBΗ`���e�p<,H9rwM^ 0�L@V	B s�R�S��R��.c���.�>�<������>�@�\� lV Xv�c�P�1�_�X�C�'Q�v	 ��O�V�������.��� O�����^ET������V��;����LPX@tƖ"O��6I�A)�<T.^�<�S��x$J-92	�ـaG�Su=w
�����x3�[W�~�h��i��Ԁ�/ ��VQ�>��Y �u�!�P��HG�cX̀=��g�SNHs+H��V�p+�*�BD����r�� 0MP�@PR��Xu/�n�-��ܳ �� ����o�c���a��B�t tN��`�&�$q��2�?1g-6]�*q9*1W���2eO,t� :�2��-1� ��$k� �gu�qP, n�����U� ���X��WC�tK��S���+��>$��x,&0tS��Zg�A:��zӡ 0(i�>�H��L������D����A�q � ������E�>`-s9{䭆�M�Xm��VWw���x��<E�=���t  ?�^�@�~
u	SP����u@@����9u�V�F
< �N�FEA��V:cJ��&H�)+�Bt.�t �)�W��0�1�9+� 0q�U�����tH��� �:)[��� u!C�� t��Lɫ� p?�'�8��t�9�tY�� ��R \���u ǋ#��^�� SQd8wc�̀�96y�KX[� �g  �[�ø. 8x�^�� ��1��25�?�\f 誰�&%q��Y3���&©,
�7�:�W��X����X��$#! EW��d� �u|�A��I�zzFe�=A-VW��`��D ���D+�*�޾p�q�X���	_*��zS��"��C;ð$t\��@�?Lu� C���3�M* ��.H���Ft5��b�8��|6�	B�\ t�����*����DaP��)'Qb�q�An\�z)z��w��A�������0 c� ;�u���*(3��d�;�q��r	� �������� �	�L�`�R2�J3%�+Ck6�@�|�*)�A).�;ѱe�+��Ԁ�QW�ʋӋ؅H��a
�)�xɋ��/�u��`;Wu��Y�$@�@�P�F�5�[G(» K��8>$�t�q �YQ��i����NS�+�Y0�ˋ�K3��"Q�h�P�e3��{�� a����}DY�-߀���� X��65��
�6;m�,8�6��O�e`@ y
P�����X�� ��S�w�� -[�W�wY�J��w�j��B�^n�`��	Xp�ha�$�?i�8:���-ʥ�˵�������� ��p�@x~����H\ X
��P��X"Xɫ*�ț���e�
- 6_�x�� '�r�
H#��L��M�p5
,�F�E�z�23��D��å�t3D�/;E��� N��9�m���t��� �0t�V�G��F� ��C @u"���#���&9���J�83�W�6� , u~������B$��1~Guu��!�Vk�u����g��Ė[���v�����(����T���d���[ɟ��m9 T����r�(TF�Xd���PD�n#eTp��;�
�y�>$q]���E��!���i��� �mX�NF �l2V����p+�e5�y ��"A���T^� ����RQ�R�u�   ɋ>O����+�> .��NN����Z���G�a!� |� ��-+ҹ, ��L���>Rv���� ��O��%��t �L��+��V�F� 	 �u����
YH$t�Y �Q��p$�t��t�� �%���YI�ы�GQ�n�G�(l�F���y�$�$� �Ὁ6��N��m�#�	���˪���D*k�m����v0�s��؋�[�W����Q�X+�H,	d�)���@�5�'��y��Ͽ�U� ������P�.���O	p�?&�>� 6\tA1 u:(`��/�0{>&>B��{�j�Y���Q#�G��G� _��~VWL�U��vd ���6,3��묹��S�H����D�����t'pu��� �@@���k%�8���Ct�HK�N���  ��HtI��W�P%=� 7��� ���Ń�
;ir�x ���+It+���i���n�������X��3�&�mp&G�'\���XP�D���$�$���P�stA-m�zA����A,���\�t�u�u�*@%�+�Dð��W�VQ 9��� �J;�u��;�v����� _�<+�S+ws�VCqi�p�t��5�����+�]^;�r��Vk�v_}�[`��W����]�LZR �K&9t&���u�H�KIKד��V���" �aZ=� t�=v�=X��=E�+�=$ uIdA���#�;�$��X"��aC�k,�F��vZ\p��mp��;V�|Y�� ��w�Zq ��q��� �Rq�$6� S �!t
 e
y#��CC�b�L(VFFV�q0�x
,+�%�{��|Ont�Vmp����û(n8^ˡ���H釻�t=u�R��5   4 # � D  � �  c     ! ��   g     p	 W�ƴ���kn� �u `��v	XAA�����Ü�_��6x�)����d�CsH��ko�>�	�/�� t(�0��&
�S�0 ���.o�q��y[�>��*`������P ��YX��C^�VWX>2V��ot�@@�ZC)�9��@P0`7X��ƫG �u��O��	�̉%�8_a��?$�`�t�G�PP"��CS�~��XXd���9���sW�qo!����ƚ�7+ۚ�n�5^_Ą�)p
�\*��* xr��s�
�?@at,�-�.:3�4�{ �| ��ʋ6J T-NN���1�Br��-c9�y^$S���S�F
�q)[QR�$<�[6Hm/�;���"F;E�;Vqw��;v����]!'`^�3Y$�u��  ̋.q��� +�+X-��e�p��t�;<�1!�C��>�:`-s!<N����6-1'���i7u:8�9���u��R-^nTgڵA�W�f�ڀ��;�u+����Z[;�v����� \���-�Zq������;60ʶ-ur��~ ���uph tk|`��� �7uG������
 ������t43���6��30:��l��p&Tc�T��� 
�Y-�x�X
�>su�G"t˸�����<�rH�r�.�Ԭs��p
�6r��'�� ��<t2<w� ���1<w����<w�,�[��	V�6T���g��(��.]�0���n t��|��-Hvn4r�����ƨ�h��P"�rayHvn>t,rpp�9�lG�;¸�5�p��S�_��Wqc�	Ѝt0c���<u�'�X�m���
�:��-Rq"	�ptE�@"�Dr�Xqd"'u�5�2��vV�MFN����o��x��d
�!U �V� X"���1 W�����s�_��� Э����$�� w��&Ju�����>��:"Wo��-G�.q�t@.zu*���G%ڰ�.��F�y.�� ��;��6�t��d�l��P� ��H%{o�o5+�s�ԓ��]���.�� �8 % <u�@$�� ��W�d*u�'z��ge,t>(���Ȝ�6���1�fv.�GG�a����I�hs�іl_3�$�j�^����t%c�}^E*i��J�I	�(jL���)��P\@���Ó��һ�Vf.nP"�ކ�[��w�S %w�;�u;Fr�;� ���u+�'���Q3�W�Y���T�.��S	�62���� %`x;�r�;9r�+��GG�M�= �k��� ��#�YZ� N�t@�V��6D����=	 v< ������,���HH�.;K	`8�6�u�< � 6p�= r=�u�� ��;�wË�JJV=�Rr� u�6�!���r�w� �i�;6Vr��i���*z�Ē���j�;�zt�*��������+�Y�N�S���%%���/!���� �P��m��Z��9 w���5��@S���sA����x�w���I�tw��kDG�A

�)V�cQ�)�N�Ha���;�s�������靏Y��H�;�HC�!�~w[�PI��F���H9IK#[�u#�m\�p;GwG &��EuVQ�i�+�m"I��|6VV��<&9D��*4���O��Ft	Z�KL*R =ׇ���7 � � Nx2?��(V�#U�3�V��t�W[ :P��t`b�J-PW�3PbP��ˋĔ�s� Q:�t+�! 
�t�r�" ;��ß�m���)+�/�]��'���*�q�F�H�V�<~ .���r� �x	�v��V��:���%�	8�;��A����<s!��p�X����0f�V<u@	 �<s�T;�v�8�>hs\)�~�>�~� �o�#m`�W�	��X�S ��c.����INp�lYS	yR3� k�|�]!�����9o�������t%�P�r�n��F5V��3�^*46u����@�>rx������W��` tR�9+v;�r ����v��V�R��S��Z;ǋ�&�s�	C
��t
���M�0^����r�q����Jg��+�t/v ���W�Dt���!�@WT�tW����7�u��}`r��z�Ju�xR�����6mP�Pa[�5 �/. �#�  H���f�t4rUxj9�g>�72�:� ������tFP�_����t2�6p &��U"�3p9���t�����S�XX7�q���r��6 ��u�B�\���~+�  �;�v;\t�@C<" v"�GB���^R�%��q��Z �J+������t�  <w�u�t3<t�<
�t0<	uƀ> u��  �p�R���� ��+�Z�� T9Vv	����n7uJ]�N�fr�@8���V�EQP�Wr��l6�D�P��+�	W�4�W���;1H8ʠ@�@�G9<s�<+����c��oэ� ���+��6��u4�i,�	��op���H/�'`߀h����� �Z�r+�� \T�@tVHuS��'��W��G�O�D0�D�ry���%��
V]��Y8<t+����>n�t��6�����u:29F�
@0;�HHt�u��$��2xtV��X�W辀�u<;| 0O�=.u��EMA K �  G���a}踆R�ҡ��ZPVPٖHc�P*���� ��& 
�� y�����a�Ë�c,�$Q@���0"�⏤Z
����\��@�H��O����΃P*����p�b�t
�( $7 u0n�L�����Om���d��r�K�!��9���9~h�uS�Q� ��;r��뀊���闢e�� ����q襅�� ^p-;�v�<�{Ɠ^{��H�!�@{�v vq{t0�=��s	+���أ�^��l%�I�0���hf u4� �W�K4�K�5Hj� ��GrI�LZa$K��z I�V�*X kN��P��,�^��I4Q��6%��uS��z��X.h�	���!�u@� ���u8 �|� ���P��v�<�u�|4 ��6������� �uۻ�&%�<�$�u7]��L
2_+�*������#G���H�� �@�-/ Y�,ᚰeD%&�Tv�!1 j�^�۰G��}�p�������#=^\�@u
�]�����-��H�Ń>[ M�Z�����P���}L0�ia�U�+�(��(�R��ד�q

+Px�Xt��QZRq�o��ވ�X�"qx��C�p�<��ٺRS�Y��Y��<ޮ"���X�tE�>�� xN��s�M�� ���s���� ��w�7W�}~�i���xv�2�d ��� u{D�8a�v *���,q��.q��1����*q䅑$��i`-t+�>�=�+9>uTf����X �N����tvR�-u� �	;��u5�@2'���&�I�;�!�r�6�" �wgu"��)��VRW��0ve[�=\�����u���WE��������@u��9H���p3��G`� ��g��щ` ������3�QP BV��YX�3���/�t0�J������E��Q�5�p��O�1�=Q�1�}��B哰n�[���Y��M�7@T�v��f�^����\%79�����������.v&&q�F�� p�TBt7J�D�|���D ?u$��;�0�r��v��+ 6����
��PKD������<��B��l
�< u
��-v��+ϐU�N��i�C�� 1���"tLW�j�j�p;FsB�v77�vR�NX���i�*%7-Q���V�<�[w5��v�+�����?w0��!$i���u��>�adW&v�\<ey�t�����%��Ot�V��J#�w%pw�� D����Ӡhs< rJ�Z-<rB\- �<<~%|�4�n��)�O�����X��<	wt����	<w�r��0<��&q��nt< �u����E�Y���
�Ƌ�RG��V�0U��W��᪌�)n]WQ� �VW��+���r@u#d��'��>�.8���C�������sL�W���Y���7�v��z�Br2�r�F��"�����2�({���}�I:
��`�t�~�����\#���-Xf$
<
 )�tO��Pu����H��S��w������i5�C�:4T��s�"V��Y	f��)� i� �������IY*�͙@�� �6r��}��&q��  ��s�l%���z6زCr�h�lj������5���ԩz� `��t �*����+>7�y�����W#[�����|P237$���&�� u�\:�^�;�^� ����X�&	U����ΑB��cN���f���Q�q�C
聝y���5b$��%�--�[�t�F�t+rx:|��u���� �.�3^&�&��{-��;�;6�s���3����5�ȼI�tV�;�P��kS%���B�,#@Yyt�G�� wP�����b
l�1~7�M�	��!�:~@T�� w'��c���M���䒾�P3ۮFF[�Vq&�t	n�Q�T5Y,p-��*�H/YZ,�in��	��q��r�
�D�P�P���rf+UҡU=��r��6� ��Bt���W�	96.q�����_ơ��Z�s>W�*PH�sf�v�_jE���yp��� ���W������ ��n�x�^��V
^u/�J-nt(+X����.k�����6�� �_:�<5��# ��`tC6�v nJ���;�s����{�Ų�X�����,(aP����C �Z�6nb��W�[b�'� ���� r�@�܉f` �����Q���_^����� ~�$�F� t���| �v�����j�,`u�����"q$q$��aea�@�v�3��N��hu���'��c^- �Y���. Y(� ��t	���sx���.��)��Q#���U��X�EuQ�� 7Y�GY@� I6�N�;�t +�^R[&�@�%� uKKu�s7��ḥ �V������P�*���l�e�񜥢�r���u��σ�=���osqH
�M�+p�̰��[b�pn��\��t��" �����b�[���3���ΉO�8�,�i�l�~��lf;-�)��n ��萕����V��h��ħ6rd
�.82�W�!Yt\E�$Q��<�8#  f��Fu��@�t&�-�v
�F�<W6�~d�A
Pz$e�����]��n�'���I��ZLPt�W�^�(���s"�6��O����
��VS)��	��
�uOV� � ��;~�s,n��\-��	Z	�r��C
��W0���3ξ'�JV�aZ��"׸-�=*�����0W�E�NH�@D��S��@>P�s��>�]|x� <
��r�t*ҁ0:����w� ���g��=��������u��y_#����[J��`J磗�Zd�P�� �t�OFF� ����լ��S�*�I�$h+Ɉ �wO
�u ��$�*�WPRyP�H��c�+��+K�%
�u0\�W�fR�Y�W��R�WW-F�  \�-�W�o��;�xx0����*�������6����W��]d� K���Q��6�]������=��bȢe���ז���ڡ1����x���H |���������FtGN���>P��	t�	��ˢ- h'$��t ;�BuYr�+vQ���Yr>�МPE��X, =�<|=�L*�Wb�r��'I�����>Z-����C��Pf�y��#�3��
 �8����
�N�3��~���a�)��l>v ������	�Ⱥ-@\�W ���=׷�����B�  �u�5k`�=}�\-�a-%�0@u\4);xp�t�"�
��p��-�� uWP�
�\�3��	07�ǈB�-�C�k���s�v�֏�������N���C���o��3�Zx�ƽ�ky@��*��+ɋFCt"��K��O��O�K&��{���?I VW��p�61ؤ6>0���+������#�n]_�ϸ�A��� � t1�=	�V��-N.�� F���+��OO F�NN���H�VB|i�z�N����\V��������+���Z)VN�~�H��Ժ  O��,wA�6�P83��u,{���#�b��lP��pA�3 'uA�#*� ��S9����
0W�3��BW����tn�����v �%W�Xv��+���&��u
���F
��䘼"Q%s�r�����n	�v���Zvl	َ�������y���m��t"����;-���&� +�+��j�����b�ᖡ]��f��+�J�6r�����&�!�n xs�? u�,�C���n+nv�x���J�t�&
�u7���#GG�2 듗0P�{�*�e���� *�*�*܀� ��� 0	K���X+���Sb��z����� �(  ����#�a�V�@ 9��0<Fe�PW�.��s�I�#@�;�����tX[ c_6�tI�nৣ��^t>$�Ww���3u6��qha,Ͻ3��A�eW��3�+�\ؓ
�b�X/�� �J X"��� ܈9�$�W������� �P����V:  r��YX���� ��ԗ_t�Xa-�Ju@���;*q��V3� �V�P�B����t��&�����G 8t����RG+��2�"��������0�eE�� I�t �M� �.q����n���D�����������;4B��x�Ġ��P� ��Z������� ���ǦGOtD�2�{�pb���85����,�$ík�� 0�D��\�[��"u���M>![vCa����C���~Њ��%B�I�6�\���ӽ��y�ӣo���p7��t".�t=$��tnS�T[M�[��P �^ðE�r�����~ �u�V�#j�wB�	�0Y����p�v��^���2kE�3�u5���� #D]�����a��,��$	�fL��VWb�=�W�\����
���dQ�-���B.8.��  �uu�ލ��������|����ue�O����te�J*a���Q���K�*~�c��0S�  �΀qF� q��G�#p��0˚�J��H$�vt��ɨ�_��$��<����
������!���)�� YH?8n> �B���m��0�Y�6$�Rz�����D� �)�(�u��書ՙ�-���� ���� m�fE�E���m�@���t<3�u��`DW���!vm���� ���}�Y� �����W���+�� _����Ŝv�L����fH��^�M��.>VL���F��ڋ��W��;��r;���&�&)�#����/�C� Y"n��Ζ� �V-�ָTX>sRiX���p��c"���5�E�Ռ�=^r��g�i�����)  ��Q��JJ��=1�|�3$t�D*(��s@?��@�<}PSS��|�ð =�� �F�x�@��w#���?���	���	Vc	���	T	���꼊	����謝�:��MV�\)���ۋEV�>��G�܍D��Q�� < Wv,*����/hO�q�v���%�i�C_���<�?L����D��f
�NN��
�#����� 3��t"���P�d>�xR*�oNN<�HܖW�xd��3�;Ƹ� u]N�w�1R��Z24 �
��� �7����� �^��pp� t+���,%g�PVr ��d�<?3ɇN����!Q�P��S�!�j�	˗�9C���&?�O �x���T��S���@�G[��"I\�z��f߀���81'����u�t�6-� �R���ɻd�J������LûteBA�ͻ�]˩H�&�����2��H.Tu>&�$��T�A'�m��S�y��C�����̚8h�~追4�>}zHz���`E�@W�HL3���ö
.�#�A� u˄{����N6��2f��#_���T�AV�7<��-u+���% 0H�V
;�t	wV	��vP�z�+F��a}I�(�)��h�se)��%=o*�r��̉^���$� �󪉝ZTp=�~�k* ���&��&���/� �3{�  ��s�G���
 ��t�2���;�9�����ONC� ie+�+Ҭ:t:. F� G��X���0��t
���kUPI �tH�x��QΎl����B6F �d���V�6X-�p�;�s	;�s
�4���2��`V&�8$uKK�:��������t���- W�^�V��w�p��N���ƽ�p�$Z��u���9����>�-;t8m:ˡX�.�H�X@2h�s��@\����^�ڡ����S`B����[�8�t���'��u��z�H�O�ֻx�t������`�M�S���y��t 1��E�^��$�G��6S8MI����	XV�v��F���c��F��F�0�9�A��@_wGP�6��3B�
9΀n�tV���k��!�x�Ww ���z��z��t)�S�
�t����v��u� ����(t!7�ʘ)NA���G�%i����/��t&W��= �	
R$q���띆�qTyytg7����n��9�r�� �wr?VuFF��eC�Ix*d@�����  t�H�����p)��b+�u�^��D��r��a�^�pg�������5�� 	
���t��s�D�`Ƹ������1�)B
����sM�0�:)%���ƚ��;��w6��t��[���H��t���2��u�΍�@P$@���ɖ�t�M � 	 ,�-�L�t �;�v6���At!@u?�"�r�  �t��*��D� �D������� ��حҍ�[YJ�|E �.P\
��W6��! v;j>�L �+�|
��3���r�3�V�a<��w?_��R�s+�4�tU��w<rw!�~ ��P IS�FF` 葯[�A茯@$�L��œ�Q�<���Dl�AO"��֟&�QS � uSW�� ��[Y��.�S�%�0)�)���,Q��(��Y��7^&8��#1Ú�f�� K�d�z���c �N�̓�|���֜ \�^
�G�"u  �-�XV���3�3�����&�:t$߀u	C��P���^����c��F8��V� @*�O����Pu��0��\/ud���rl/����$*Q��� ���c�ۍ4c��g�)�.�371�6��`X"�&��Ö�~&�&�ˋ��(�qm� ��-��F�Q��+�r�L� �Z )�% @��	  ����X2�f y\�3F���6��Ҋ�.�.V�F� �"��%+ ���"0 1C t4+��"�� F� �t�(8F�wu&���YՈ�6,F�����:���ו�u8X���?r	?�`������������!��,��^�Z[���� ��q�*��>j+����pj����'	)ݸ��ހ�M�KX"������g�謤V>e�/g	L�S	��N �:	��!(�əf�p���~�}#���n�����zr���x��r�n������3#�"[B��,@@g�/sHH1����Y�n��6� ��ez+ r���Ǉ�,����|�'|��z�v���}�v2��2u���,������	�E��E�R�a�D��a��&.^��#�i�����88��I�d�� @��f+��� >,\$�$P�f�G�=�t^�g+�1����.l��GƆ�Z��2�9��sH���*�\��s�b��.45�ǿ5�G�.N8'�r���jh k�> t%~��o�2�
�<���>�� 
� CA<6�\OG=�Nn��~8�G
�W	�0u��D��H <��F�F�*�8v]�>Fx,
�>}�F�%�tEM r��vr-�\bw&i
Si��bF'"��F�j k��F�$s����8�A����\=��-�7h���t<`�13��J� ���H���̳�?�N������7�(ʹ�	�M��VVE����t<�K�ƛp�/R�X�-0b��-�W8X踘�b��t+��Zt�>���oft�;V`�B2d	��n`;ď�&�q����
*4��n��Z�H��&� #(��j�� ���3ێ��&�ܬ8� t� �&����gǏ�8 ��(�j��1|���×5`d��5�56�Gy͘��u%7��KG���1��n�$?� ���CC��s�.��0t!��'�7t���HtHв����;�\��\�3�at�2�c\H; �qK�f�:0��>q�?q O���6��q<�]�)�8�WߗE�n�u&:� ��r�4���H��- � o��6tWN��M\�D� F��A�N�� �lz5t����p���h<�u44�z����h-� ˰=�ۘh���N�6�%/ ��A���V�31	f:�t�e�*��"ڸ� <�zn�u�[3��\���<�	����x3X�YB�����k���t�n���RHFw_^�B���H&u������u�H#�f���PSQR2�m 3�"�.ZY[RX���f�3����S�_2�3Ɂ>D4vI3� lJ������#������������ �����0���$�&>�'��[�&	�� �@Us�y$����#ы�����a9V�S�WD>`���N)�I*�a�D+�?0�:�1�5:�07�+9�,�e�F30~a<��|kܝ$�{��F�a�[�,�6�h �ds�����w�q�P�'��b�`s���$�>�t����$'E�_�,�����E P �P��'�.�T���1;�p u�E�ƼǏ]>�>�l��pj�G�S"��F�K(:�m}2�=GN���G���
3�F��%~�t�*%!&�$���~�u�bu(�g��v�������,7� /� �/�F���.xF��l��eOM뼊I#,[3�L4!D�iF��<	1y{F�D?3o%3uSL�~� SC*��)��uP�p�p�R��f$��^��7C�u8z��*ˠ.P���:r)�o��	*�`w&2��.�j(?	i�V�� �W��F�2T����$��3$�
OH&!1 �X#@k��Lu���8�R$'��X��!cG �wR(�."�J�)�o��7xBd���u�2��h��!���Gp w��7�2��/��S<cu'�&�C)t09�*t	tt�n
t
�ӏ3`C
'u1�<�B
9r v.a�Vt)Wt$��=��= r
�\vv���Od�wGͥ` ���[!�{;E~w�������&������ˢ`��;Z-Z=W@Xx��83C�U�{�#�I'o@r�gHM
'��			�jR		�	��	�V��
�^� g|@C�@(�A@s � Y5=�%����� D�����J0�q�����=m������3��E5�� 3C��6��	:	3��	17�@Z �@�������ay)E��uW �����5��LC�{@;�u@`���o"
���U�aH��W�W�׼�&�Mn'F��>|��آ�E�4�J�03��)$�*#3N*|I���J�2&	2��qU�� ��n�0� d� �55� ������ 5J3�� <�33�����3 ���
�  �s�&/Ϫ8
��\fkxR�~(���u���<��� 6�� �����> X����� Z�rx�4S >�%+17�=ǧ ɒ ��,I�OGW���~<�%w�F�\j	��m�v��*�P�P� �W�ϋF= .� =s=T=tp=(���!�S�<
�B~`)������f�a0�c��t$��~
�
��v�j��\�F
;
�Hr�v�#�X��a���$ �
R�' /G�sd����)�6-0�:I�	�""�

��=���{t�=	�=
a�=�����@?

� ����m��t�^F��h-2���q�00Z]�Đ  � � �G�=��8��$a��p�H�i*��0,�&VSQ�0J;�yd{�� {�2���� 5���	�f����54��;#�^һc ;u�y��p;+�;Oa� C+W;Gs�v�7V�E^u#�s�f�bhT�<j���t���S�)��;u�*���0�*�0���,\�p&+�[9�.�N��-A1�3��H�>�R���q�!�a��� 
Ht�6�p����v�% Vl��R�
T�<9�V��]jE^��U���^�mO�O<�O�#�Cu�b�����L�F���@[};>VquH8t��+�WV�譧
���9tț,w
8+89�qc+��i��p�X���2��du��G�����&��ta�P�tP���P� F;�Üd- �A

�+�P��PS��*��@P�~�$�Z-H;�t	� ������"V���q�X.�����u��
Er��3�_�%
��b��j�C�tK���Y�7���2�����4�oVW={Qq#Q�rx;�GEt���O ���lSP�0�7��u�o:�n���t�+��z�6b�dG�@vH�;�tP���6` ���q�s���I�p�+��J���	=HP�j�x�Bt+b���;0�B��7B/���/AtGBuJX��0聤<��ހ>�t)��p##�i�e����v�ftN!x��_��!똚�ma~3� �O�[ �*q'H�E�5+и S � ̏�U�
�m���)�� \����f�����X�>W��PDx���tȡD�X ��w6��rjg� �_8�G�yݠ��A�+��H�Po�A�Pq ,�ȡ^�u}wdΩ���S�x��%�,�z��2���Q�M
$t�-���-�e���\Ct4KݘvRqV� TZq����J c-P���X��ۆ (�%߀<i<K��ˊ��-�^ +��~�0z�xc;�v*WWr�mr�G
7KA�P��w���D�Y��������2��� �#�B��'������ _<�! � `�FE
r�{$�^�L�H����E'B� ���lǇ�O�=�3�"0�0PM���
eW��� �(�6&��u+  ۊ#��.��X������� ���� F!d��)� �]9Yt�n9�
�e\�>Z��Xq��@lf���M�Vq���b5�qm!�� �ut1�p�@�a��/���.3�)�^=I�U����8�=&LU� l��8��<r�yn�L5w&�r'D�R�8!�/
!�VȀ���W��X��#��"���9uR9��	l�2e�L���`�+��#�fƬ�Q�P^�Y��
��"i�I�ǖ�V�"��$6�-�"��q�3�>ͷ��w�T�z"�BMVP~g�V��u"g�!7�L��	"�n��B��V�;ӳ��Ӈ3)R��dV݈�@���
�u	|\�9�/Lo���]D	��  +������N�Q�i��&ndsBNVW�4�4t���� �O*O	'� �A
�H��&`\� >���6Z�>-Nx	;�)���F�\F+VE�TX�^5P
 vP�J�S `�]�ON*�M�sMF�wA<豫��1+�@R�S���#���tN���w��m耺 #�3�&���`�j�V����%�����ΐt �O�c�c�X��+� F�L�D�v^!t�VW�B��u��� = �t+�D�|3�d�VQ�QSR�<t?�I�g���~��+a ��R�4s}cf ��\�L����3IVh_5;�����/:9G� �?z �W�������"٢���)R3���n�-Z&�V�*!W�������NӸ ���^�2@Z��v���|o�Ϧ����t�������$�M<�����sJZ,�z�CDpQy���rQ2��te��kD�	����~5��.�+�~��P���$r�{br�(�	Xr������/(���~��\Q��,��+�=�5�Ԙ!����eb!���(���j3Ġ���pK��zԦ̀�#�
 �(9�k��$_���d�#�_����ꌐe����*��z�F���˶���1��	t�Fdt�ÐWwB�>�6��}9~u�^��_�O$�$�7��
�D*�D	t���t2v2��+��2m�2*�.*��y&Ru&�v�u�$�-WD���Ӊ��E�G���T*�m����#�pF�X�G2\��G8���HǸ �6�T
	)�	A
y�r��#^�z��*�d�"���\�����i.piHP�����+�	������&�PH0��=..Y>�W�/l/HH�W1l1��l1�������E<�0:� ����*�+ȃ�QTc�,Q���U�a��#�TPM���S�>���mʜ�}uC`��4�i<��I=-��4��Q	z��� Y�A� �~�ٛ�x	��X:�jz�=����B|�}�!V5㐝��@��	�)	'T��@��0#W�SS����� �� O	� [�F��<rZztT�w�3tj�[	�A�2�Gǂ`��������&gbLr@�D��`J_�_K	m�MA~�M���[*Y���B$%���B��Vh��iR�!&������"" �'F� 	p ��j��B^�B)�Dx�RV�R�u
m��I@;�q�����oΨ8���: R9�t+����̉	�>(�1��`R �d ���L����0�	h^�	�R^(��V�C�W �2l��$���G$0
*G�G�80G	�%Y4$���(�F���8�����V�:�/����%�N�$Q���f P�q 
 ��%�$n�Qlȫ^��\�Db� �uu2.0_��x��<*�!�7�>
?
=
.�:*��@]-;�>��c�wuQv��W�E�f�E�E�E�B�N���2��@�*�^�0!�G��~�;hSH����Q���Ci�>�(+�u:Ƌ ��F��N�� W����`��u1�ml�N��P3�F�- ;$G!���A;GN9Ar�u�<w	�!P���=^� ���}��������'��'��"���@*��"�A�6��i� Rh�n ���Ղ
�~	�gV��4�63�2�J��O?Q�y�������������LU�
m0*
���|�l��W? ��+���$H~D�OVfm�&4�VA �G����V���H��w���
讅���%2��p�<3������F�6�]��LL	RG`V���'�9J�H^�\�W��(k ��V�. ��9F
t!;$������$���$�8l�l"�9ud� w�~ u�L�e��M��"s�VHP0M���AɊ�,��	��bes�C]G
��4��S�_����̡u'p� Nt�,���D����
�� ��Pܔ���ķ�	 Ý���v��q�$yt
��0<���9!t�&+]� ���op3F�hSV�oI�S�P�&�U�K��J�=�h�Q|h}hl����2k)1�h�	�}c9u�F�P&d��d�;�RTQ��,��'8���d=���@�o�O��6�������I9s�@����&dǆ��! �@��㉿B*Wb�u�>b.�u���J*�I`b{'�+��^˹����*\�v4qQR"��G�^���\kO��@�||㬫-]JY�N�:���~���b/�N�"p��y�yB� �+
I��"�EoN���6���\H�,�"0�8Fs�)
V$&���g�w� ���Q5�v�X*/^����N��@���Ut9��=\�^�G�i�B��r��\�R�������������'"���'�Ճ| u��������
���_^H���F��D�w���M�8�8'�!8U��-ہ� L}��x�+�V��qQM9���c9$@�	��[��>�r0y��>G;`�
�S�uW��Q�
W?��uYY�W��6�F�p�߹��v=I(=S�&===	de��Q�aî�K��p�º�l�?�>48�F
`u2�&�Q96t#�$Z� ����-��`���m���Q*��²;^�B��~u%
@��E�`M��� ���Y�y9sƼu!�����^�G��?S1u�7�o8U�~^%I�E�F�[QU�yYhF�f?,zhe1�y�7�d��#Ai��Agf��c����1�|]*�G� ��� �GΊN*�;��u�%u
���>�^�&,�6�8ܯB��N	�f�O�)� Rƀ�2��P����m�f�6x���ITW�-4p�%�~Lń >N ���I�1��I���r�,/I�DI���^ � �̶�
��|�t����l�����Y@ ���QuS;�7�\v!m�p�Yp��@�N� u��QeE �
��W$G��
g�bs��mׇ�̬ �a�Uh�e蠫�,t�
��aM4nj�j� =� ��t�9rD@˶��1N|�C E���/���4yI�1	�'�8�t�K*,�L*�з�:�K,T�0���-#,�㈚��($������%#�[W ׌A	V��H0���낄���"�m���C���d�BXLq}P�Z#�@��?�u��pI-�W�N��7����E|0�
 ��+v����D������� �P�� ����� !)���\��u�qJ���tt�A����-H)f����o�.��c��v�n��tmr��v[k�y����
���tw����?Ks�@+����#g�h��SV�IN��)��,O;	 �?�F�@x;Ā�T�p��Ub@���� ��7�1b�D$��"�� ��s�8���8`��.28r��DFV�z�����������,����=N2� "����]��EWV	N��
�:R^s>vz��f��� $�� ��F����LX"���S��}kExbKM	0��^@�?��1���C9���NN�'X$[#�H���N�1 �F����
�� �+ҹ �
 ���0�O�=�6�Q�R�:��/�/)W//��/u>�Lu� R%PF�P��r�#�P�*'���5��V0���=����"D F� |2�bV�kY� a}�D������p��k�� ���
+�R ��^s�P +� }Vz���"͵>'�����s���Y?Ð�5��0J�F�(�0W�C�20&JP4H)<���y�O$>�7?\�W����;tF��N���>��%��O��}
��	B" �^����}���P,�� ��c(�%���ۯOz;Qb�C��+�V� prn����O��㻚��n�NWS�d�� �^R�H
 �u�\��w
��[_� 3�8&|uH}��H{ˢ�^�r �s�X4/�nx����O�\�2��v�0��9����>�-3}V��w@C |H�̀��xt;X��p	���5�-���!��8s���Ĵ���� ׈�#�Qn6 W&F�� �q�-�;�w��%4i��@�S��l��a��W���.y�m;���L�e�X����pP�u1�4��`$����5H���w�{1�����]T�J�f[���y��
=�(�{��M ;�v��z��-�Zqf�QT�Vq4Xq��o;�.�*�ye�>>��l��=�����1���� �W���u+��B� +ɊIx7t5� 1X����(lR��H
4����;�9av�����  ��_���uKxS�:ph�p��˚�o��������}+VII��Ps=0�XP���>���zC +ЉV��^�S�H>^�VS-�[��;�r��:��&C��aj�+��E����K�W�� x� �� ��� �t����P��0�+�v^�rQ�R�6"VPWH��_Y�C2� �7x<t<$t��	�� 6G�_+���=������ t@IQ�SY3�á�U�? HE���S���+��.�Y�[�����O������u ��-
�t���-t@g� � H�.���I
���.������r
�x�_'�;ـ#rX7tP�&a8��oS�q�^�[� !�@�GX�Os;�����-u���qd��@��!~��� ��Xt����+bDn�"c���f���Oy�ff?���j�����O�J�2n@뱚J�� ��R��ݍF�P��K`���Q7��`���#1L�d%q'7N�۸��*���utJ�(�6��/�r��wO͆������{�(��6s�Pb�H��rN�Q�R�}C}1/0~�#�j6����v�'*J�P:G"���>N�U=��)�
|�Q+����eH)��|�P5|��4�c� 
`Fu=�  �N<R$T �ٗ�6�=#j�2�>�5�5O�[�EU�|GM4�����~6F�%F�N�o؋�O����!9�S��uHd�>4x��|Ϡ.��"q	d16=�M'�z��^�&��|�5D�Ś8h��$�&r��<�s�44z����w������p��u$u �#tu_��t4��&��Ү{ ����I&*Xs�užZ��-�iRp�A�2�1��U����a3�-� �yn)y�		�		=V��_/�I*V����b2P��^����p�JNVW��z @u� ��`� �����FH�$P��� �-"�V��Nvp/�N�F������IƘ1p� yZۻ�l��h=R `S��NZ�@*��RV��jZ T�� *Ӌ��
�L��:�SR�D�"q&�v����4 u��NG0sW�ρ��5�	�ƪ�_GX0��#�-%v� -��t*�:�v ����ي����*�*ڀa<���	�.>���c�PQRW���\`��uF.l����  v
�|:uFFKK_ZNYX�?a\�@��-ۡ��x*�  ���������u�@	���X�3�k� Ѣ&~1E��'1РC�H���d$�&K�q" � 1����I�ފ�	�V�I��8����� u�G��I��Ɨ#@�{�Wqx��A��k���N�)���?\u�� G ;�s[W�0�OoE\
�u��kW�%z�I����&~-԰ r���K_�pKu�tu�2H��TA��|'o�m�m;'�b�� �*H���� p� ��'P�.����qn4Aqvxq�����
r��|5+B-��L13��1mz�1�t#&6�(�T��H/�a�$�h���N׌j��G�8�"x���0��ƒ�S9�-s���6TsRs�g��@����d$b�{P�Ů�����tQ�-�������m���Gh��W0����0�R�Ƹv`�&�b.aKs ��q��ƺ�{���/��t׿IaJj]��q9!s#�p����t��$�T/�
�/l�FL
��&
�fKY�1��7��-�: ��եL���0��� ��;Ek���v���LZ��R���W�P#`��q��6Wv-�~q�e�e���D$< D��ى��K�Ø/���˫��ٸg36�tN�<A����E;�xg���'����!콨w�`���`,~�u��?�F�PK֎����X&���1~
��t2��Hp1q��!����>��Mt��W��=��o!
� f�x�e�P�S6� ��;��݁�����0��>HDBA��; �R-�9�����bB	�A�����2�G �
�<,�.��t辬�Ӹ���-�����D}�g��"@~P�M�"�[�H/E.��B#R��wġwꁹ����6P����{����7��4X���
�{�8��\8��1BҚb��X"�Dj�b&b������O@�!N��%LJ����T��^�d�j�޽t%�
�h ���(��8�p2��r�ƃ�N��P���L�}u<��f� H=t2O��t�%����&je��J�y�AA�jҧ=$no-^t���3��WP{b�  e������� 4�d�:p�$�>n����C�^
�^��jj�q��u����� ,)�u0�q8�Du���:�Z��dF�O*����Č$�=�3$� ��(v�M�����J��О����_�Q��G���x��T�4 rA�9!��0+DT��w�&�v��"�m�;� Q��ƃ��:�!�-�������6�����<����d��X��\���V�[3��u�O�A�q��f�`ё�#uʙ�'�
�9S�GYj���J7�_&PZsA[��#�!{�U��'��}�7ɇ�ƚ ���6"����~�YJ	-3�1W�ɡ�9QR��:W����Q��C7��b$�\���������pGr#U�z5�Ϟ� ��
� ߢ^���|� �A��%!4�dnF0�cG��9�r�Q;3M��kP�F��w�\w��J�������2�@-d-4	�>�4���BR�E�o�3$�wN�T]g̶���$E�!N���A �	ϒ�AV�����C��Q=�� =�w<�[�w	����`��W��-��-��I�%��Zs���'��{�!�2�SgQhuQ�t����� �h�7���q�37��B��\^��T	�m��
�A����{'�]:�%����(�Lg/]���VV'B=m�xL�;=��t��� �{I+�u�>��	6�:�A�D3͙Vy��5�����uH���=	z&�0t!=&=(�O1'�_	�@� Q@��FXY�Y��#��������-j����������M$EoD��E�eJ�1E͸	@#�����_�I�6!"�q�g��X��w��a B�ː�!sdNø ==�<3���7��JT#�3���f��PSQRM�i͵=
��
�1#ZY[X>T�<�>�1 3VW�N�V�@1@��_^6�m?�{�6�?�vV׿�V�E}$V&A�U�[S�� �[ ��L� �x +�P���[L�� �,	p	� �`3���� �}[��SPVS�z� �ng�=B�QB�B=uT�8�D=`tS;��=��=P �u7�5V�M�.  �k^���t�P��� .�����&	�}-|�c��	F�=��/G	����X�#�=�l }4���W�؎��>Ȋ��Oj_�˾'L�*�� �D��X�]��D	���MP5SQ��
�
��SQ��Y��ø� �PIWPS��J�>��� ;VWS�0�![<rV�  � 3�� �3��u��  ����'�Ϭ�<\tw</uw�
� {��t"����	��0�`t�<S����[��9��s�  "T-�L~6{;���Ma(a����P�D�w�D�
P��{�.�P��?�2���~)�)%��$��d��#��
#�>t��q�Z�u
�����$��Tp/��P�QB�E 8�W�}�  ū����&	����  �<	�^�*MV�@�^�' XPoVL$� �GL�Z������x�~�"���D$�nq& Ս|(�V�6���q�  �.GN$��j�z� �u��:��!��t��eI�- 	� u�y�NL��T���:��cs� p"{v�'Pקg���5�IO�!-�fp��^%�@�9�����ff9�"Fr�Z���������9��u��r�Y?u��en��[��Ä%On�S���zZ)�鲬J�� l�[� )h��u���|J�i�"�8%�dw��O{ �C�I�x� �lt��g��ƃ"4�OpO�Z^y) J�F� ~]���0O�ZF�QQ�PwS>��;��;�>$q:�:��.�)���-3a���-+��g��;Y!3Dz?���'� �b0	��
H��t@],�p~r��I�!G�ZPq�Z�˙r>1�ę�4JP�����)��r�m��VIr����)���C�x���%���)X�G�F�B��F�n�\/�%�]� h�� �V�����6ck�C�K�6������uU���Md�uL���[ B����"\���fG�y/ <�	��~�y�t;�W���0�)��7ն!�~v^`���������j��C���2�"9�2u&.u) 	R	����)t�\C���w���  ?�v�%�<-u���D8F|�j����l�t�%�֛^�� ��	��PW�2��
Y�	�,�A\�*2V��E��T*R��/�.�Fԣ����� ����U2v9�j9�� ����-�v�v�G X� ��[�Ф���F:� 3+][!*�PPPyd�����yc븋6�BӘ�B�dN,"��B�HTt)�H�)�	E��` ��쳸*P�F��D�f�B�2,�3��0���Z-HH�Ш�Nr��r�|1k����ĳ���VW��U�Ƣ!�rU�$@��N�>'	  ~ �2���р�B����/p"	�^��8	C��	(	*�чo�6�YWW�V(+�X����h�E>�N*�,P*��TG�rڸ�.h(����@3!'	�
�����yI++�KO���~��Q��]��^erĳ����3+wIG��������O�+�R�+�]؉���;�*
�����W��@�� �D��5��2���/��2 #]�f��_�_�}��<�N��������甕����1���1�_�Ո:��j����l?v��v#Ĵ&I�*�#���4V�8����ɿ%4�&���� �Bc���b4�4��ib�+BB^�NBRBTB��BBV:�BXB�J�/���J� �q�7CQD
�
�$O�6�x����E��2&)�j�G@�T@��A��Ү�{^�A�=d5=� UI����ӗ�s8(���n�pn�~@j�r��T�W�l`����Ȓ���P�R�2��t%�Զ��;Htm�[���b���-n����tu������P��cw���� Jj����M���Z9 ��pԽ�S�6�T���!%m�K�o]68��^b!4�i<�8a:f@��wf%�\;\�v�}���R�1B����U11�1�Ͳ � $��Y��SSPãQ��X
�bP��������r��.�5��]�.��E$.�������A�� �8�|�Ȃ�-u�z vz�x��.���_�� tw:Hg�VbX���|� d:� �>�a`s to�>8th��P�.CQ!
'� �
���+�� n�~
'r'�w@���lwI)��-UdI����;�ջ�4?Z���L�G1L�(��P��j
'�{��.t�c�(�I3�~���
��� �� ��0 SG�_ ��������`E�9�
t��ϣH��������"n_��_�O�Q^�^���$a7	������W��! �
�>�q��#�b ��++���#��0�#� 3�8�=�	'	� ���@�P�> Pո����衦���:�k�HWV�X�����m��� ���� �2���^�6�,�,��)&� *� ���+�����y+}�3<$t8pr�3W�Y���6G�1d�8�DIK�rsḮ�T���3�V���P�������G(����k9&J�X9��w�y?sM��c"�h��egv�T��1$"�&ѵ5�r^Ъ&(/� #�'�+���& �,��ށ��S������NI��)Q�׆�ظ�Zy`��aF�z�n4�A.6���*����'��y�Lŝ 	Y� ���d��G
JԿE*�`�y�8�y��d(�����iY��  �a��Wg@2go���3�t_���d�
�x�e�xuk�cH���8Bu���*�1�;��f�����-^橲}A�����C���Lq���.Xw��cݩق�x�u�Nn���u���~7����W��7��n�!!��p�' ��+J*t�!Q ��� ��Г���(�bO���~�;I���	�UT>;S[t<���s�d�)lRed��"��XvE$�$�t$�	���4bs9XsCV�6��K$蘦 L�w �tG�a�rq' �eYQ����r9F���Z^6�6tq� ^֩=����0·�wA��<�L�����8�@p�
�j �Ӵ�*	�xa�O��V2^�$�^�g��@��V�LL3F���e�I��B��:o�ͱd"U �y��{u�-
�m73B�Q~�-�g  +�^�&*G�ȈF��׆A:s����!�G�Ǹw�R���K�
����|��	p#b��@Uu�`*n�bd��Une��VSä�)��%� =jm	�R�H� � 8�In+� �	�8'P=����3ȭ����.�+^�dkP!?(^:7��� t�g ,�#I��8!(Z*G(*�Z0�s���^�6�H�Z��#�Y�����&�n`!��bs�E'T��yy ���8�#�0j��8=`��៺;{	���4�Pk��Vk�%�<`��������)*���|l�@�;��`*�\���@jH�v������P+S,t)�u�� �U	Vw�	u�T	��Ur_���P������;F*�tF�� �9YV��t�!�+A�����!D��m?h�Lr0@�ÚX2��T��ȃ�2Q-��yU�W��=�;�L=� �&EWb�� �(4��CUvM�囄��@o��fJ�*��]H�ZwS��Wt6�s*���)��aC���)����wQ��������M�nI`*���������\���m���*U���ؐ<㓓��l����{x����y�ϭ6p_�	�wBC 88X;5ATU�n�a�|����e���4{n
2�ք*W`����F��~~
+vFS�K�$�~V���ɚR�윋�� �&h��+F"�4�F��9��w�Z>�/v/���;�Ԧ/�t�E��&9m���u �>6��w4=��� [GN�z���. ��a�HF>HG�؀?:uQ(��N�V�g$���!)H�Rt`�9v�rv3m��j/�k��(D���'�"�y�<:t)�)��������0�^f
�B�iL덺�©� S�� �P1�u(�s=��	;�=G���M�
�+�[�
㍌�r���C�tS���(��$��<D�1�v�z�2�WzUP�*G��  F.1Ț^���F,73�0=h��  ^4�x�#ֹ#��*\���O	*���7���C W�;�������hZb��X^������� �@�W <�s"P%�   ����.�X$����@�3����#Ó>3AV���l�W��E?^A����x�F.���lg��.�I>` ) ��!A2�L�n����D�:\4$�,0@�дG#�*�� DU�sHZ  �VRR�: Z��߀�A�+g*��p(qS����@ &��Z�;Z-JF�+�.<�u��m���ĊĢ��uD`Z��w6T�� p&�:�t*R�	 �P� XP��T� ����Z&�*�~�q�Er�ش>��x�~��E�� u��v XPP��R0C�N�&
&�
 "
 ��U��E��A  ��A��A��A��C��E�0 �E��EcI��I��I�  �A��O��O��O��U��  U�YY��O��A��I��O  ��U��N�AA�OO��A�#�O��P��Y� `Vo��[o�aA��^�AarF
�x�*�<Xs%�� ��n.��C:�t�:�9�.�G�L�=���	%�P���D�����3�8$+O���3�øi��V0��5��
O��
��M� w������ qV��P��6V�[2VSS} -gP|x�d�H'�6� p�	藬�D��x�����b�b�e�iT ��4H�P��#���;��g�IXJk2F�G�Mt��Kz����a   á@t'% � � <
t�F Ht�D�	�G�9 �@�����$m��W����p3��򯷻 S��=3�_`�V���,#�B��t��%��W��S�@%���[�PV���=���ڑq��u�G�>���+ΉL2��qJ�$c�P��F2�SQ�ܙ��Z2�V����3L���5	�Y���P�	X���� Mɖ�G'@_^$1�C:���q@�f(���d(3��6��\�����6ǀeSPw�:[Y�����G���D;!u>; D#|8�h(;�w1M  ����8��w����[��F1������Y�듡p6H�l�	KQ��!�_辛���LO�s�������t�09�u�t���q9��!��*�y<t	 ���R��ִ�N�a��v�Yc��Al��}����wZ������u~`t!R<(#&U��t�JbN���P�.5P�/��A[B|<$O�ՑS[tRGD'Ë�<��toLe
��)���u`/^��u6nE�M��:W��	G �.W�
�?\쿓{� 8��f������KXu
�G �x���.��j_��/c
D�k���Uu�-�A��) �!u"��	PR�x@7ZYJS��	[
)PB�Oà�V��r�x��A�1���"�u�.�Q�4 up"�FV��^AW0 �����%$<t
3�8R��"!Ab,��_A��QVWS����Ρ@u�vS��Gp� ���L<4�� ���#Q3��6*�S8<R���?��S�@t#H�  �s�"#>�!�ǂ�J���L�Xg���:�). ���:r�r�  q�s5s!s�s�s+tht�A�t`�%ӋN ��؁���s&DVM �.���t� =�֊ǘ �q2��qS-�V�pP�+��= ��` ��j=
��0Q�p���r=�d �=uI��	u=�F���Hs1��J�`��ް뙀t!
�u	 r�}�k�.�; \�;F
u���nm�ƍ�P��+&��Z�n���^� X EDIT.HLP HE
�	QBASIC�V�Z-�, t�Ͼ�!lJ��'Sp�K���t�������^�#1�[�"S��P����D!;���"!��荽X� �NA�f�\(d(&��3���EI��$�9u�u	��[�-��p��5`W�68j(������73�8!B0�À>�' uX���td��Z��7� Ii_ �rW_�S��W�ORPP�� [W.(���i���l$BM�~����WV�b������u@�9� t-�;ۋg%��@H'�^�HU��$u����C�B�Ir٘��o8��A=�b�h�A)��x�ty��e�b�U�\@P�9X�����,�� ��% #S�D�on�� ���|���W3  ɊG�2�C;u;aW%� �� ����r��l�� N$��w2�2�afpZX2E>�xՉ=���3��X �P� �<�	 *S�*E��S��[t�(4[4Fd#8Ou��j[�A��_�1�@���3�qPSM��� RQ�}�7���f(��y@-6HP8-]��JH��* Eu:�s3ґ��W�0 8	P���Y7n; �� �u)�6�q�~�
��/�W�@��[��C��K;^� v1����"5<X�_^F��}�j�*�C�HQjjt	V^�G[�j�_ 6Q�m�G�;f&��s�aP3�;�F���f�� �(��<:u
 �:fuۋ�FF=,X�X?8A0�Y?�G��P�P�]VRU��u�(q�H�����'$��	�â:R 	O[;�u�x���J�)3�h  �^���-�F`E!u��8*:�>H`xץ�`tI� ���tC� 9#<<����3��a�5�+���$�kPH蒲��9O2��J ����! �� 9G���Ý+��H���rn%΁k�7 ��z���X��� ,%�.�*�6E;A!�t �D ��q����Is�<`�l�#O���~$t�.C(Ɖ�(�lOu��B+ H�DtG��(�T��\�B�  1��3�&�&�Gp� W	�6 ��q�>Ap�/R�^_�3[ 	W�F��0��u���u��
|@
� v����P�̀?kފ�����u=Q�i /�u+=
 s&I<.1E� t@F�B6BF	p�B�)��	��W�p!<dY$�F��D���uò�2 T�|�|�|�|  �|�|}}EJ &+'/009+�9`% 1'])_*8^9F  DD	J]#_$�2^3@I2_r^+�3� ���c��w!���.���|.�  ��F.�:�r:�r��@C ����ή���|�V.*2�$�U���X��R��'0�!� ȃ?t� ��OQ����Tr� ��[�D�u�(03���-=�}�P]��?�&S�9&� �V��W�6�衜_���<!N�t�������Z���8�Ra F��&B ��%/��v~70�ڒ�;F���д=�!s�e�q�^�-���.6~�8~�hL݂�$4~A�)�&���<$t�1v��9�x�]�*3� ���A��I`VQ��u���"�+��t3Y.�R�f6^)�GG� �u�i@��L��W��0a�����_I0R���P��7P��>�X[[	����G�%Š/G\���g���#a��NSX0W�F=Sֶ�A�!['���x �aOW��F����5�~�� �R��������iK�u�%
V�Rj��WV�=�((�7����-}Pz�B� (�p/SVP��,��vL�P�����d$|8�}E�$W@��O [�Ă[�T$�@��%��,u�S�E�,9��'t�^6��
^��.�y��'��i�C�VA4v�� y<I¾d(�&W�&w@��� @"�>pW��g(t��O�5� �֏_�=�y���0&�s�p�'��5�[�CİL i��er��p��c�[����X�%cVf!�p��C��L#�5��&��� 9A3������� ��Î���&�5GG���'���8�����(+�Y���La���wڥ �z�����Pc���Z�Z؃�y�S�g �J�����`�Y��s�
�Ld�[�V�};P-`G� � nr;]�V
ͷw�~�|�}��+،"��+����������<�J��NO���F��G�Ə�I�d����6?�~�%d�l{�� 7�ʋ�%?�N p�3�RRQ����y��@ �0��� �3ɇ�cQ���脙^�{B���?���}6> �,Btl�J��V���`��/�D�X'��,��8Q <	� B�!Yr`��V�?s��@���K��Rf�>�u���		�3r�s�=#�Pm ������&��  ��J�� 0 =XR��.��[�����yL��Ơ8��ZX�p�WV��t@ �+�����狅4�� ��؊�6������7�F��|�
`!�v�,�w��-,��HdHf�HgHH�>jwD+̂D6t:��")R���"$|�+��d2ː�
��GH�C��  ��. ���	3Y�a"<^6�Fv��	�9	r%vD���T()F䀴�H���� 3�T+PPg-�EnIW�L>
v*�^
g�W8� ;W rw;G
vS*�B�A�ؙ� 5������8ډV�m��9�vUSR� �P��$��n��σ^� h�����n�n�w�n�A��1ȋ�9�N�����#����:0i4�u�����G�|�Ki�i��E��(D����~�P��� �f� r$�S�� ��?��Z�E�ESb?"�*b�&5 &�&�����y2vo�V�F
X �)9SE��q�
�F�����;�vl?�
�Kp�&V���!\o�^e�_����@7@�!�g����Rj��a(�0� ����r�����g*L��v�cĉX@+�5���1��VK��tJ��̞����K�^!y�&�e�9�$�	�/7���s D�G0�F�ot���y�"^=K��
���ib��<���&f	\@U(�j����F���k
�
(�M�1�����sQ�� 8�+��ډN��^�ㄶ�SQ8����)�'0@iDH�-�^�9�m+ܽ�9Fr{�$�@�uS�w�P$;�x��Z�n��s�J�N���n�HcJ� ˂��$��i���9� x��UV�"�K+��b�X��nb��l��,�2�2�)>yL)d�{U�I�V�F� ^A�~
u�<� �����f*���d*��~�|�?�� �Q4 �������CY&�\ 
#I��GI?|A+���	���GżV^;G<�,��7���h�
��  �Y�+P�!	�%��La�*E�)1��V�9wr9's䍈��x--���� ���O�wG )�N��v�V��Q蟢�i�8�!V���/�����^���NcT�������yu�:�9"OR����{]�zt-�zP��t*r*���2�$������n��p*���EE�l  �2t�~��B��EJu���I_:S�V  �[�BEGHMNQR +� (� Y�<{a�o$<ar>	=���  �6� �65�� �^�  3Ҭ<	t�< t�r4</t3�iuE��N�v����^�F3�G# r+���# 1w�6�?����1�$_� �� 0u	���.�� �`Lh 8u�iq��D
�r��~��}���� ��
X@;�v�~x�x�� y vk/u��Y��%__=BFu��� ��&�� %�OHu��!�<Iu���0CDu6�&`��=UNu���YY��I��x��C.:u&C'/��N�y���OR ����N�=DCu�OMu�14��HEu�L<�Pu�
��N�d�t_� x�2t =u�
M��v���0��&
�� ��¾�  I�? X"�X3$�ɺ�6�
��e4� �� ��.�g.������M�P�"5��n�2	D�o ��q�������� ؎��^�����^�K��  �C+ދ˃�(|�' ��&�6�   ��-�/ � PQ��PS�������-Pj�Rt�X�� �L���$#C� #�_�/��`�	&��/���/$q5S�t0 ��-+�ø ��K��
�g����J{�c@(��H�XRVW������u\�<+]G��;�y�s"�a�gSٚ�Y �rY[Z��pt��X��_^��u��T��*R ��t.KK������u ;Ws�4r[��= wwQVઋw�-^Yù�:p[�># `�������f�*�����=  �����o�V�$�=�vԇ�AA�7r!��c=)]n�ati27\u^�� �WYZ�s�J�\ݷ�i7����KP���Ӈ9V�L55,��Q��GA��0%�Dp]�1��m� �&k=3�\A�|s�
��v%p�At`w� ^�@E 6P;Ev&VP�+�s#�P�u(����Y�]�0R^[����ʩX � ��$�!�u� \r���AN�_|Mq��,�B��8�n�U6&�eI�W	�":�g7�N�� 4�+N��k���c��g��-+]�6~D8)�F=..�)���h.�>�C�}B�RL�3_Oș8� �3ҋ߉��Gvs�v���u�P)������RcP�[���~� �t
S��[��
��0���b5+������ ^�5B�v]��~ ;�sB� =��G=�~xi� t7( � u r�a �'$� ";�v��軽���A-���_�&��Ef��%P+� �s��[�r�5WP��鍀 ��<X��;���S��g�Q��ێ�n������ @U��M
RF8)��+��1��AT�06�_���$OzCh��
�l���� 4 
�t'���u2� �� ��Z ;�s
���V

��N +H"��P �7ږ�Pá fq�d��-�`�lfb���@��6�8h ��B��lJ��
 t= �u=��-���� ��1F3Ɉ6�-��: ��`թ- t�b�+��Ή`�-S�3�Z�>vt�%��`�x 4u3#tӋ>� `->�-�}�u9�6���6�K,��F;�w
�{K����D���L��a���`��[hR�w�� �]�u���������g�V��jq  ��E6�-}�E�	�JPnC؂)Re�BX"�F|-�� ``G���&�q���\.����Qw �y���+?s��Os�O,����j1�"���^�v=h��u��� ~�����QA�|B���"�H��9n�
;�60<�OR�I�T�f�� �����SW���c .�_[�u���v� #�  �� P�2҈)� 3驩����� �&$� ¨�Ǽ��z|���P����`�a�R z&P|*��y��������t��\���M � 3� sG�h�B���<�N�6�0�R�#)Z�fY[X��p�(� a�Dr�$  #+�tF�>
#;>#t �}�=uE��=  {����������6/"#��l0�
5��* �D�#_^XË;6F�<t:2�+tF�D�D+���W
\��94�+�9�1�(+})l~���XK�I�Du? ���t+�=�4��+���D�QW=Eph��G3���
0D�_Y��\'��'�Q��L���L�����pi 9&ZBb�Q��/��T"'����+�p��F �L�cNO�+56FG�	��t	�}w�iV�B;�����^_z;�08<�\+�&;`p!&�|� \*\�G��`�0�Y �T w�wV�7DCC��^�>�BA�׸\�u	k�vt�,؞��+ك���10��5��Ot��04s:`
��p�W6؋ȇa�vA�O�5�?f���9��_��'RW�����I�Dd�r�
���-|����u�U�ܐ �l�����OO������
3���@*�E� _�����S��"���&��ݙ�u�Ha�3�4N
rPW\9E|�)�_N�9Ӌu: l�E�;
�h#t��xj� �t����F�|��  �4��K�o �#y��#��q	�P� C��
�`fó��ff	
ffffff(23ff4567ff89:;ff=>?@ffCDEFffGHIJfvKL�oݐ�1�D*#D�����y��  ���u��� �T�=��#�:�1Lc�3�]H땳�
0�t�"%����΃>;9�"t�XZ� Ai��Î�2���ټ �# F���Ӌ�;)u�O���������S�
S�(�� 8� �`=` X"[�>�t�vB�ld�`��[SS�,#,G  ����S���� X� �f��P�>S�6
 ���OB;���ڬ��� ��^�R�д�!Zû&;���N��0Y����X�	V����������PS w���	��������b�D�s %���s�G�#�,1��=��QSRQ,S�  �N���r7���^V6 �#��s�i(喍� [YZ#A	�\�LԠ�[�s�j�#[���V耱]�lF�:S� �W�����	 %���� ȋ	�w����� ��P��e P�L��4s0$��� Q4r$PVS����[^X$�(`IV�^�5� f��w�w�[SQ?̸�>����r:  A�b������7;�w,��	��~
#��E�Rb�" �Z�t'Qu3 �+�r,W�[ o7
�E�p�����gO0�K+�4����_������ ���������|���7��ח���D��-k�[�<7V��t� ��;�r#+�F��InN�O�`X�BMȉ�;��%�>'� s�#�#��+��B�9#uA�?�X��� ������+7r8  P4r.�6P�J X� s�@( ar���N�N �x[��R l��� X���:C��?� |�@<D@9��jV�A;�rD;�9�v���<F� ���.; �����r )t3�� ���x�t
;�#6�I^������`% ��ƽ-��4n`I @�r����QWR�=�;t0���� �>��Z_Y� x�|�G;�t/(� �>�P�L��+��+���
W���20�N�� ���O��+ϋ�L@MÊ��_���t����a��RSVl;9��v���$ �^[Z�WD����r;�rt�Z�("��2�_����  ���Ë�3ɋ����0 ��/��������|]�@�� ��V�d��\�^$���s8��L�uS �h� ���;:3�&8�t�0 Kw�	 &�2��� WQSP�� ����X[Y_]�*�q n&:�8 �56�}���,�u  ��G	@u�G��������6;r]w"����K>\�t��X����&(w0!rE&NN�  �� KK;�vݖ^+@D��D�u	������PVCt  ���# sGBP�.g��s�(pH���(2�'"#��t)= �t$;�w t�C+�X����s��f���)��`5$#�;K #����`;	w5�&W"@t �-���H���	A�]����[�!M�����5D�h��;�vʋ�E�:r{���b���k���u���;���uG7=��h,W�&�"���"%�Ǘ�A���{@ ���+�tN�L5�>c�'�W�PV�`;�tr' ���� ��+�H`84�s��H�9S�3 �;�rFguvg�	��(�+<]
v)���.��؉�+p��I�f'[��e~x8}��@� �� {��+�>7b&�+VS6���\�����w��\_��T ��^úRL�T�!a\�3�9(t��)9u���X��V�7 �_밁��sNXAw� �; �� �������H�6 @Q��V���q�W����A��M?�=�89G|X�� �)Mr�sʨ�s��9��Ç���$WX�$����ʋ���!�O��jX�����WQN�xf" �?�17q6�&;���r#$#wDP ��A�ɀ��L�;�t�|������ �R�Q3�B��JYS���� �F��@t�;M�L8���Y�B�;�@�t$����uǕ
��Aa����HZ�O�<s�#�t�����u��� s���\�]`��;�	��;s�-]z!��[����r���+�t�����q� �X&#���^$�v���%�����E�#J��;؜tK�J"�V&I˳tCtD8����2;�w.p0�� *r�0��"��7
�s:�C_ӦF�6��I ���d��3���@�M��V����`�z^�$���V�F�*,#��dr`�� `�|u	�PP��� ��.#^��6 86� �4�6(�p#�*#�� ��} ��%��� � ��=
r�4Ԉ�0�7��:P�Xt)�a�.	� �7!���ub�5G�U��>�CrR���602Y�Z�t�O� ���_�ɨ���%���k��~l�U�!+����^�#�]ˋ  ��Q�Y����Z ��L��p�Wԧ*-�� t&�ź��  ;�v&;Os	S| [�N�>� ��:_��Qd�Y+��\_�3��W}OH1�,�>�7�%
��� �G��Fg,�r��������j��)�\�0���E�T�8�u9�t�z���s�� � �ܚ*����À4u��~>� �� 1��@@;�r�˝9�fF�
  \�� % ��0<����
,�#��#��	�0���'�'���A $�;�r�4�K � û����Bá���P�Ja�s��أ������� ����(��ɛ5�(���2�nf(��V
n� ��&�1��ڻ.��E��r�16/,�Vp ���X6�>> �44U>Y->"a��p�{X3���<�D�.�M :V�`sB u�����3�����68���P@P���(  ��W� ��t&�	�x& �s&V�v�Pl��^_���5F0"�)�M�Hs
l��4>�)�I:
oQ V��2�d&!>-�R��n�v��$����E`�|��
 ��G���P�gBx�h� �&�� �8��9 ���x���3F&�;t$t���9�h&��u�h�60��ډ�BD� &X� �64�J&3�܈c&b&�o�3�3�@t�t&�� ��=R��x�&�� � � ���| Z;�s�H
�t	���1 U���r&�p&�f�&%u���=��	��6�R��� �� ��+k#��x!+��i#x���o�=	+m`�#�����Z� Q�J}Yt
�yr�T��� �rG��G>X"� �8@���؜���&h��&�P�r�����D/�pD� :����8[�  ��ʡd&��� ���t���`��i3��6G 2�+ƣn&WV� ;1 ^_;�s��.�a�N� G��%��9k  �sz�p�>j&�l&J  k����m.j�ڦ� zu�߇։�&�6��+���3f�ѣ=+E�~����ƴ���!��c=u"�>beu��UgXHt�6�q0އ>N6��a�JP��� �TQ;p&t%f�rfr8DrG D���Ԁ�!t��@u��@��t��u��n= �%��8�邐z�� 89��3�@+���2���� r�^����t���C� � r�$� d�P�60#P�#p�X+ � Z}	=��~�3 ����v���r+Z[Zf�&RSs��}�8�Ep����R ���\�Ȣ�3���VS�CtCu5p����CC;�t� $�=����v��� Ȥ�]����Ã� ^ز�� ����>��u @�W^�� #�}�-  �����VQ�U#�V�
a� '�[� `�0N����u����Y��@^������;  �s!�+��+��0�<5  r�O���<:rB���A�1�����A  *�Ԁ� �3#�jP� `  �PSRM�?5�! 0.��.��� �%Z[X�PR.��Z��İy� .��-2� 6�7�^���5� 2�t��ظX"��v#���V������7r	8lxi .�<�h.�F�P��Y����:� 7��2��ޜu����S�W�<�<� ȧ�[�� �'&�2n ��� �� ��   �� M� �� �� ��   �� �("T7"B�!N�!X ��S�"��!P�! ��^���>�ʺ�	5	�/x �)���2<+t <-��3�'3R��, t�n��3Y����u\ �� R���� 8Z3����>+�<�,y�>3&0RQ�)�XZR�-�h[[QPSE� �1I��ZN�&sA&OBP��I[���rO�������'���1�x# ð@��� ���q72���&������(�o2=6  ����a2XR�aZr,�����Sr% (2��
s0�  .4s�� s	�t���&W�{� �û  ���u���f�Ɛ��J��� �s���B�s�X ar�ɀ�sİZ��  ����1<Au���1�h�Zy�;�r�`(�����2�(g�)�!��)&�#�: �� :�1�E���1&�=�0�?�2[@c����� 6��2�ꊆ�����#� �����"R���1#.�ˁ�]�6/�>� q`'2�8����
�t^ˋ�6\�V�W�,�7:ι��s���
�a��뺹
�������tz  #^.P��gҞI��U �r�/M�%���0��ݼ�SZ����4fT���r;�oG2H�=��
���u�Ͻ%"^�� ���N�O3U
�G͍ vS3ҭ+xT@��⒭+���[��g
���.r5OtW��� �u(��r\�wG�3˲�  �B�ٌW�7w
�(�8k�%PR`l/B�wM���ZXt
�Ew��Ü����2���C� �'_^� ]�-���$�3�3N:�u�SU<����EE�����'���� '�� +G|�;}� ���� ��][#�rw$	���?�� �+��'���Ǝ��߃@ċ��`fZ]��'�U& �.��3�=�̘��V�0yE �t�*Ww������BW�GH�h�=	B%��d:O�W6�-(ωw�w �t�7P�D�Y�:�Ռ��5�.�ӝ�])�M-O?*�'n'^S?��Ga[A�FȎ��I�{���t� u�L:�6b#�w^�`)�#,� �������`4V�x�)�$r�^�3)���l�G�B�^��6�hz'!S�� V �[����s�WU �u�NPRQ�� �e��� X�8 +�5�s<&u ��e� <Ht  �<OtN����u3�+��I�UASVU���*]/;t�u��yϲ۫ ��;�t�ɀ�� �u��[���㊪at ��
`u5�\��7�S�7�9<#u�4��)<!u� ���<%u���u��,� %���,�N@ud����#�t"�
��- ��K�Vu:�D��t?jo;}�V���.>t:���0R�.07����Ztt���%����Gq�=]� �; ��<"�,N� ��3ɬ:�t
���A��,�<��u��O� :��f�A  ì��< t�<	t�<
 �t��i�Ì1���%�� a= v����ݬ� 8��r  �������R�3�+�0Z;�5�-� 0��~#�K���0�D��.�	���2#�
�� ����Itg8!��E+)��ڴ-gu�H�T�d��40����
@>00�붾ˌ_����982�=���e���=��< 90t+Б/������'x���@s�L&��P���C�^&�� �')\&,#v
M����)RP�$�v8;UrX�ጃ� X�X�:~q�r�&�l��&O��L��z4Y��o��"���rQ�`M_Y���^�r[]Ԥ����0�@"N�����^
�8e�A�{�n7�W�bS�����2��kHиQ��z)Ȫ��+��Oߨ�{�(s�[p�ZYUR����ڣU����]�� &��*n�.+�Z�Fh���]]V/;`�3ɡe#���� �i#�k#+��u#@���_�!g�D!m!o!U�w!D&I|�S�B\`&� b̦[��5\1�ג��~�ƒ,i�n�L�g�1�I�qsq�T�W�&��&�U��_��>N&���+�"�y�&U�Y�*1I�� `|]�&L�PSQ�7CQD��BYC��(5���T���L��[X�\���sҨA% � N�,��(�t�f*�46�A��#�=�BuR���#��� �� &e���� ��I��+���@9�5�gF4@���[��9P�8.%
�!�:>u
�#�#z�H#�#-��#w
�=�#�aB&�p�uPzeQTH�fmq#�L�c�HQ��s�( ��r�SQ�>� �sr7�^[h�R�	)9G	�gO�F	� �t�ñ�=�"��#XZ��G	�rH� �#��>���-��^��D�Ԑt�M௚P,�>�2ᴭ��ި�h~D�(� s���7�u3D	薏�}�H�u�苐���82���;�|��k#;mo����Ñ������z�g RP�_���\Q$�'	��Zr����&P�"N�L�T �
�#t���-����
q#
�+��I9�����3���7P^�J��� ��SR���Z[�'��'�á;�t(�֒q�9,r	�;�t���6-�99g��� �e�ˊ�^�V�� 		���e�t� �~ u��B�'k_p�n��&b@���H�L:���

HM�E''� ���t�]� ��P@�ˣ���ΣL&O"QI��RJEN���@�-%��(�a�m����$��� <�t���]����� �u9�&�&�� ,VCtKt*  x(;�w$R�:�Zw�� C3Ҋ�*Ի����d�Ӷ��Oï�Jʜ�N`NO=��!��P�/g����b��N�b�^�@.\ ��0� S�Ls���t[�*�1�t�85r��#Q��S[t#� �bt0���&�`�5��8����c����	<|ҍt���� �t<� tI�L�T	R���(�P&�J�4E��[TW��d P ��B �Y���\�k% \�����<Z	 �S����=��o���g���W]�\*��3ٹ����r��P�N��~8'����p��M��k[A)W*� �^<
w6� Hx0Y� p�*P� �S2t"d&ZPR���~��� �4���.- ����  �< s�<r�<t�<t w�<s�S� J��{?[r���A�o�Jn�t���v��������.��1Dȏ��= �111&1� <�������$��F�-$
��
#�
���T�#^��s�e�i#�
�(,e��>�&�Y�+����#n"SnIE2�\�  �� 5e3]4  �4
@3s4A3�4�  4�4�44	!3:3 M��3�J�ۉ�S'������'�� 0�� ��ێ��&�$8��%t�&��[X���Fu�1���r�����u	`<�t����u� �<u����<�t����g���b �� ��>tt跊6 u`��#�]ٲ  �@H��$ <�u̸�Ý�n<���`��� ��>�S�P����~��
��~R�R� ����t����Z�v���.�Pp/�, <� ����
����,_C�Z�̽�Gu�  �V����1���1t.8��#�����1��� .�T���^\� �a��� +˾,)����À6��ñ����6�gt�5�+��.J��g$����S����S�  t�) r!�+�#�l�~
� �r%�K ��bɌGZt��)ʁ��
����(S���A6����'~ ����[� �/���[�|7Ĉ��QY��\�S�
x+g�#��t�`&�gCOVK�*�i>!!?!$8ډ�#)I�+�1n��])pң�H� � ��Ƈ5%J^� #���� �_*%!�U�� c��<�� Ճ S�K�c��{��u�������m�p����Ss�H�#KC�H�r��C�6~� s@Չ����[�cL�c��Qxr�CJE'y'Pd  <0r<9v<Ar<Zv (<ar<zv���sru��#�b8�#��0H�+��Q�N ���R܅���<l�譒C��(\c6+ˬQ��蚒-Y�3�8.`��H�$' " �P��$<< th���u�6��J�H4E���輔:&u<
]=����
�1�	`�;\;��L�C;\�� ��L
C,���"��D
#m
+DD3�  Ë+	�9H
�c���Kr!^]X����%�[v�V]���w������������_ e��P�g�V	�	M 3�I �� �	?K  �YZ
�t
�t̊�:���v�>넽� ���r���` u�:�w�蠁�� �rG�6�R�DIu�Ί�Z� 6Cu��( 1�t1��  u'� �"K��wC�ô �<r�w�&.�� %舃r"� ��tP��X�9]h�JW���FH���Ӧ:��v�������s���?��w��c�ݛ�٢��t�hA���p�*��� 2{' �II�°F� �+ ߩQ���z����<	��� ��Y����p=���
��` �0u��#P���mX$��iN
@�
�u!JH4�s��B@ Ɋ��I�$=c� ���;X"�<��2">��;Aut��% A����
��XP��@�"�|	�&C�ӹ�R�L 1��	�V2�~�� �"��'@'���Q ������YS�[  u��G�܋��ۓ_��d 1"�^�t$�D��V�
u u> |�u89�d3t�rl���� ,f 2��� ��\ �����������drюF8����!��<" f�,u� �"z� �$:��"t!<tF<|?�'pS��� ��a���u �:�t:�w�P �ds�`�4�)/c�{'-���Gl0<�z4x�c o�I�Ҵ��c^2����7��@���*z`��_"���u���� R�@��	�T�ڋ�Z� �û;�t	VS.�����ޑRYt��� �$��_W��+E��A�����^D�%�A���Q[�ga
�] ��� $�6�#�>�#+s}��+ZG���$��0 3��^
  $�~&�H�
$GG&�l��9�#E��pe���z$p�?������S�`�&[�=�$�����:EG=8��#t; ���� ����  ����.��r�w���7v��'8�It@|��A��'�u��8�<@�n��&��6$o����Z�9 YXS�X�D���I�h�	$�Q�t�;��t ����!�c�.?�.GS����$+��e��  w�ȸTP�RP��:��
�
�a
���\]� ����M�\�N�3������!�Y�t߂�S �x�����6S�t$	 t�p'�r3�'�(Q�aY[;ȹE�d�� ������atr���[��d�F  �f��N���yD'|�\���KF&���FH&���`����*��������F �F6�+%JZg�Θ=SR��� �� >�

J&Q�7�˂v	
R�d]0 ����ZY~(�f,�QaLS2�E[yY��+�1,�<|�>}u;t���Wj��.Cw� �U��uQ�*�
7���)i#��r�&mas�� ��� �y+뽩r+���{�>�>�eWPS+ً����+� �� R���X���<����x@��Ƌ�K��@�BP�Xt;n�3�y����
���� ������u��D������� !*��
`Z����M��>���6�x����6��i��*V��# 
�VU;�~�`��+�+ӳ}{��ȋ�۳i`w���ډJ' �.<';�}#���ࣰF'+��H'�A�:'��2�9m�/\��t!0�A��(��+��)%o%
r���q5Sz�5�yM�?(�������s�e	�GI� qy��"~���]�A�_yn�H�~t)�Y�٘���&��# �L��Q ��z��@K�O�}��M  �� �B& ��~�WVQ��\#E���� � �^9�SM� ���QS�EP���r s
�c2�X[Y����^;�Z��t&�S��� �����%�Q����3��C��p��}ԋ�;��3ɒ���3�j3e��we�!r��
 �  FÜ�$�$�$0�:'M2��� ���r
����������#��t� @��ӊ�$��׊�=�Q$�s[VWU�RGf�>b�6<'Y6�aC!.HSV6 H%u^[����u�_�)]V��94k�99��`SW>w_a�>�6�>�6�?�>A'��A���.;'�� ��@'�{ ������ "c���o2��c��M�l A���<��:1�� I ����@r0~���P����Sx�X�%�%  <&�'"���s���y������2/"�0/�E�Q&&Î> ^BBBBBnBi  BsBuBzB2�����.����A���#$����
�& %G�"�&g���M%0 �$F�������v�&���u��B��"�x$<B>&	�A����*DUc�`�mb���<?_�]�
]7��]V�3�V ���5w�}�+;�r)L�AN"�F�@ �A��Wċ�1�
�x�  
�Kt&��s���0Ʊ"�TG���N��t��#O0�t
�� 5"� 5E��S�M�.GF@6;j�3�?�2�"�t	���E� �U�����;>V'tY ��r	���t*	����|*r':%�=�=s� A?.L����s.�qqJG�%l0K�D�M:.�ET'w����v�0�ݲ�1�����������Z2�]U���<��'muMt`�G��X'u�DU's�3��� A $A"$jIU�ŀ4蓊|g.0.t[w�UH�G���>�tO9�!v7h��ju�2������U*���� 7"�"�u�%%� �C&������t��`rv�0�vr�� Q�����Y��Z���Պ�*��6ˠ��V�,$x$���D ���k��s
���y%6F'kKu��> F��&2N "�&02�4�)E��&%H'>7�� ��+�s.$(� f٦ � i���i��n���ss&�7��^�Ȯ�Lȷ�}��f&@�@~@�@~�#����1�Q�����
�� _Љ<'��������������U�6L'LO�H)��NmJP:'v�)�qV� �V���7��Q>��ǓBah`^�&�,"�����*������9>Ar4�� x�޷����H ���0B�J|	`D�&�'��J�$ú��<���1>#����j  j��r���#���4F�E����t�#.J'�ǽ�!7�B �~��G"琊���/ڿ�*�/C0L���g�I��=�D���zE'�*G<�  �,G���1G.׊��A�=���4�w�ʗ�J�<b�J�<�6�RDUR��=�a�<J��L������6�&$Z�8x<[�o��Ʉ7�Ӷ�PF�=,F�7ZX�3w,�fw�@;wL<NP"�4J�hX2����W���JB��!
� �x2�
�Kt)��p�ĥ�&�GQh3��Ą��u��\ '�-��;G У�P 3����D)��b(�hU ��D W  VS� � 2�Ѝ&$��8%O�G�	O���
��*$4Ny��[^p��� P'�V'R'���X'�PW��Ћ��>KZw��O��F�C>_X�R`��A���@�2��!3�Z"�&0ĻD�	��(�Q:��u9yƃ�i��Z&�
��M��!��'�'�]'	���@  �=�� �t.G
 �OO���͊î', euLV�\�1��S��=B`� �qc��~@�e%K��s�ť���U[+  FW�`m���G���_�������"B����Ջ���;0�=���Ý��u
�u �B��s�����"��B��+G�!��%%�Wr%�%2�0�"�u�tF�5W� Ou�"�2�t��0ȀU���0:'S�>2$�<��u:� xgt#F� �/�3�":�� *$uE��s�� $u�[
�St��F�7�Ʊ���[�я19]ZjD�(t���N�N��������KW;�$N*4�� QW�M�&��u�N�0���� ��2�s�P��RJ8JX�(�O���.������b�/*3�2/x`�/�`m��D�vF�&�OI�
F�>��5= G G �������^��� ;6VY�$	�2	��� ���ͽ��U�*�U#2��w	vLu�&%<���uH���OE#��Gt���k����}�2�VEtM� �;����:W��8i��U��4� ^_
�t	2���R�����5b7�#�7�Y`hXJU�C�^�Jt`��㵀��8���qR�6̤B'VjDu��3��+��8�t &���E8(OuMT�\��� ��_WV�����0������� ������Zx�6�q�o�  � �89:;<=>?yO�O(�Z' `�F$W�61 � �Z�U��(����0= ���;�t�?r�4�� (����: 0'w�
�
�u�:(��:u
�"�V��2�'W����)A;�r���̐��V�	���C_
3�QbYr'�)P�*��NN�Kzo,,S!= �![r��$�Y�_�-�w@3��䴥`u�+$s�$��,M )Nk�)��)Ɯ)���`*�z6H�&
咡P�'�+�R�a+�6� ��诵���> t�Ӌ;��u�R�f���I�;#XHx��t
u�?	 �G�l���w��۶.���3��D �[� ���s^J�

  �uC��Q[�ڋ_�O `�^S����+G���- UP���[����Ě#���D}6#=b]�9�t�u�ǀ%���]�3ɉ1�e�+��X�P� s��Hx+_�	�/ +P���L���`V��'�T�<Bu>��q<Iu7� �<Nu0�=�+^�L ��d�X� ��������a��v��^�[�\Xi w^�i����<��Wì�	���<"\o
�0��qvR�P?@L>Q�Q R����<�u� �� ÈT������S`���ĘH��z��4)Xn��>��V ��� �� ��D)��&.���P{�l���`��h�a R������ u�2��_���� �%SP�� ��`�[�0���D��!Ǯ��^�p�A �uᦛ!;�ضv'u�E�����e��t��MB��< �|��@P�
�g�ֺ:�r �< r��{l_����@� 8}%��Ŋ�Md���wL�K�㊇Y�@r��M����6u� ��X �N�0�P����W�0GPVW��� <�����X���_^� H߃���	�ÐF�_[�≶@��V���QJJ)�C�
^�{W�O 02�3����gdx`�Ƌ�	r�r	�Q����_����G� ��t8��RP�7u3���u��<�% SP��/�X  Z+��r^[Y+�ʇ�6ʓr]�R�5a�3۹ x ������ �9&��S�[���� �>7f'���
���tE0��ȋ).�t70~:�tC����s ��QCw�,�s� s%ܟ� �? M�.�g��ٷ��d��� �[e*�6;'2im������m*����O+�5&<��3ҋ��ˣ�&�[!�t��S�7��0�w���R�<	t��
l[�m���  5���<=tJ<+t�<- wu���������g�  p��<;t�<9w�?�Ë����,0���8����t����� ���V����� A�^Â�?	s�ݖr�Z�	���W���.�~�]?<[�O� �T�r;�s��8�P#�򘑀�V�u��m�ڿ� �ο�o��� w��OI|>h ��|7�~�V  ��};�s$�+��p�;�r�^
;v	�wG��a��6��<����;�m�	5��@yÚ�=X"�.��2���s�`���Sk .��9�����" [��P��a ˶ �ʱ[�r��
������r�C"FH�Ý�3�� ���&u��:�H� ����swQV �<���^Y��Zr��`�P���.�<u?08��x0 �{�P�tS�   ^�@�� ��
�&��F��&	 W�/��$?��&���&�䢗	���&��sIYr�0���	]��9�]� t��Ǳ�Ӱ�DE����~�;4�B
S���`g��6]8�!���~&�| ���6�&+tCr��]N<I�;� ,�R�5 �΁���}`���N�΃W��>�ke �3���&��t�FS�a5[��0��1��r�3�r�T�6[�>� cۊ��5��0��|���u�'�2~2A��,e�p�K
�u<J  D�&Q��YQ�� ��  2���U����Y��&�8�H��<As����&��H���%�E�鸳MJ���:/v�x�]��(T\�����r�[��v�&݁>t PR���X2���+�s�ڈ�/8Pq���ZXڞ(# &Y6�7 �}��;�w��>LPta�����VE /��2�uq� ��!Ku��#/�sF?Q�]uW~�k���
�u7��ˈ
i9��*x�(��u��22�:(v2�7�4V� j��~9���12���:>*w����}[:���FG���7H�'I#�u�SR���K���p�5O=	�-��H&�I�b���= 
0�8���&��D  ���&��&Z[�8zRV��1	� 9sԡ\@� #��X����>�P�\;UXf�b���TPt!�q .?U���������P������Љ6]HQ ���^�UӋ^�Ȅ �g)�7��5�ʒ�<�� �
�XZ���}t d��� �r$��Ƽ�JJ
�%��5�^9�P�� D�PQ����>d/ s4&��'���� HC�h����r�X* >���b��y�����i��YZB��S�Q�$���s ��*��]W�S���&�[�,���2�|S%��
"Ft��ؼ�_Xx�x�tC�}P�D^�fC!*!Wr�!"�<b�,B$���..�v��m��(�\����&��!���0���0�h�� �k<u��a ZuKtW��� u/�@�� �ϰr[�l#�� Ha�HL'tN�,�qj�g�? MFHH�Ԁ� ΀�(X$�΋/-��"Gj..GLK5�=�h�n	�k@ud�5 ����*̑���P �Yr��n��YZ[�����[�t[[RQ˒!fv�t!:��~���^F\**�r:�s	f�û�����w�p�W�̓�<D3D�*"?y��@��Z)�9 `ܾ�tY�x VW�>Z$OO����
� �� B����_^�8��O���c����-�� !e9�~Q�'W �A��  �^Yupug�� ZP�w�u�X�y� O@��^$�b$S���� �`tG�J [�=@�\$�u���t1��H�]� �� �ы+�3	��Rn��Y�h��	��v�����xJ��6 aP b+����U�6�3���$�:ot��" ���5����I�"�"���  JË�� �<\t�C<  ��+�΋��\�� �7���� ��"!�  ��<#t@<&t�It�<+ ��t�D�<.tE<_t�E�:u�<y<*u ��� F��r�u�I��Fb6Fǳ @SS8��P�<,���@��(#���l��(�$/$ x �N�<^^u#�| RrH���������uFI�_$�Z��u���:-�t�wZU�I����s\��6^$�鏬���P�+�4���vP�0~���\�X$,]yD�� ;�<]��O �% ��+��� ����ۉV� 3���tC�>�2#�	�+�u��u7�ߋ���|�����3�a#����  �0u������  �M� �Z�]$*�<�� u��y,���:���@b�@nA�� E*ǀ� �F��Ǌ����B@ �;H������0�t�%G�*i��v<v�V�o��(��%�m� ��
��������� �&#�� t���*�	���<t  �$�����|��u�0 ����u�,��0���x����
I�xx�.�t_~( l�����
�~�&��]t<P�E+  :uH�^� p�y�۴-���d�v�.t�?������
00�1~��%�X�o�㞪� �3#�+ƠwH����
u��.b �2Ȭ� �+2�I��N���a�`H�  ���-�� `:�=�y0�Ԁ�  2�-;9�*�%8}6 �W`��j)�ᗋڡ��ء&�A	>n)2���dx<�!_�7s�@�46r)��5��=ty��3��G��X �}�Jb�� ���9�P��3�6)[�$��W ���a��OO;� ������򮒯w���_�=���"�� S5�@`Y��r�~���$?0ZM�4P�v
'XF��ef%q66ds�����C [SVŎ�M ���t*N ���[+���+8p��R �Ϯ,�t��M ȧ�ը�̨=�;�U���$6֋u� dS�s3X"_6gm	W�2���^��9��`FF�/9�W�-0 ���s���Y�౪b� �" � ���vV�p��4�~��\,ǽ,+� ���3���  [X��B09��wn��7脱X�+b�?���O�k��2�H�P��^
�~��jv6 ��%j�EJy;�<�>�&uK�+ʓ��0�}~-���(�u$z� �����u�+هڄ,��Q ����3��L��d�S(��c�Ҳ0�L=��ϑ���?���O�
�K�|��lJ��|��  ��+�q���T0 �
;¥��觰�Dv�|Ju��m�;�B!,�p�!ٲ (1�t	%T| ��ˊ�蕯A���� ۫������Y������  M�S�_X�7���ZR^�������R�FN ���G���az�AlZsx��t��S��� ���u�:�r:$�4 ���[�HI��=�d_#���)��  0��tAO��+W�0t
�O��tɐI�蓯�t���V)�� �菹���d%��࿑j��Y����vAiȀXv%�v�ËN�d����Ø�+�s�	ǲ���p���SVQ��B�PW ���t�PWV�c��T�<MVrY��N�+�u�� ��F����Q�@ƀ���s�����S���ܤRXR $mZ�3�VSPR�)1n|(��g�t�\������c*%����}�[� �2f�W�	�	� e�K
���=� �8r�NwW ��B��o����=�2�׿�l��FS��W�M�!~�!a�$!\r�_��*{h�����WQ*�Fj}N����PR�QTX���W�7)�DXXs@F@�F �a>F2E�8�S�g�YS���;ðg�ٰa��~
�  h��&���CC��P���2�! ��*��tH@(� :�s �*��ߙ��#p�Ĵ ���� 3� �UtS����UP��X��aJ�'��k`#�J&�oL�i#��m#�����*r:� �uB�g)�M� s��CU����CmYQg�y_��K��`&���R��N������&��&Z��A���1Y�Zá;~�|�	&|�6~	�|
�<	'|��2�9�~6�@'}9f��~o`� u̽�1����%�'�1��2��]]˟5�]56�Ӟ�t����+�s�? ��+���KYBD �SCRN�CONS�M1x�2�LPT1��2�3�PIPE� � F�N
��\8���9�h$K�A B�A�H���  � SRV80�W��� I~��  :u�I�V�A�"�� �>f$P��J-@:���pe� tI[2�Q�FO�}�\  �\�Y�� �s���U�; �w"<.u���s�  s-��u���!� u �f�x �=�\<*t<?u&�sL+uD�2�B3$v8
	r��.�E��C���O<J�%vG�.  6C����_+ϊ�n�^|��� ��WQ�v)���t�Y_���iuOO��u��p��a�O4;�r��0\�G�� �d$� �</�W�uI� A��� w����R�_ô�!�A:�Q�^�#�Gr^Y{�� �w�?rw+�:u%����i&�tV�`���T��U^����^͕QU�Ѱ�ø��0"��k�p  �l����'m	����n$�(% ��H�����  l$�6%�R �B%���������[������kS��z-��> �t��� ���Q��Y���@��.�^����  P�ʊ���t�j$��� 3���F7 �p���S���tǜ  C p�-X"�W�G�q�N�F��:�{�}P�o���8ku.1�ɭ(0@����% �\�����
�����\�;�p^u;�sX�������L��HH�9^��9[;w'�P� ��"^�Kx �:�s��� 5�pty�V��ѭ��2�  �^Æ���� ����xt�V)+C���ƶڧ~���WdS�� ��7AxΆ��&�� }����%��:��$u\����c��T=�(P�%X$4qc�F 
R��2�S�x��[Z�0�Du��ttn�d�5Ã�tPV8����l���g�t	�n���*�2,��
�0p,r�À���v��'3H�ûn$��^g�  ֦ �<	v*@��%���   �%�/������t�$��%�.�6�`�<�t��㋟0�)u�>��[` �n�P#��tM0�� �L3ۀ>�%u{:�<K� ��4��i�%����������m��[.=��L��7Ô����PR�!� �!�S�5�!. �/8�.�:�[�o�%Z�3�-$�-X�UWV@P.�<�Mt�0d�u�y�m�"l��u�y����E����`��!���)�%Ǎ֫ �c�X^_].�.�VW{������ :����v@�׋���8���Q	� ����Y��Ѓ�&�����������=8bN�N(�+<�C�t6<�t9���S�9;1&�*�S �"�&��+ _ك� wԉ�sɈ,�v��SQ RV���%�  ��dt'���\�T ؈t�l
:�t�	�T�"��H��^ZY���� ���%nVPt �x<s���QW%.��p  _Y��X^�.q5q<q �Zq�pqypL��RP��wq�	�X�Z� ��`uǁ
 � ����C��� \��	�� ���O�%����)+�m+++����|�%��@3��@�y��n���u!S  �����t������ ����	��%��	[&F(/�/� R�����r�����)��Zc�J�w� 2 %��PSQW3  Ɏٻ�'�VI�ێ���`��%<�!��uf�%��E��o
&ED �Ğ2u��+p���@�#(�u�w$Qr-�	� �
��A��a������y��  �_Y[X!�����`n0<7uZ�P2f
x?{� uN�<Wr��tI<c X0�7�u��)�  ������dr"��%�1���u.�
SS[r

���������3n	��ÈQ<Eu	uqJF�� �6��/<Fuc�-�'�'!(�,t* ,���g[�Vk��r) F�����v� ������%������	 ����`���2������ J�����ء��`n �asu� �P�Hp��������p�l�X>����PS�3E��KyCt.! Cu�6��� l��t�����(r��
�~��u�[dA��&e�K�*�6� H�%�$ �� ���i�9&� �t��%��%�cG�&�&����0 f
����l ��:� z u� 	/���65 &�.�rXX�A�� �ُ�4�]2A�N�zH�B��>Δ�l
�tƩ��1�s �(��Z�awS��p!c���0� ��M��V�#�A���_^[��)E`�5�����O.�)���`u�����5A�BCD�EFGM  �v�au�Tu�Du�9u�)  uX�t<u>u �d��d;�qߕ��_���0����s�'�I����s=�n0sR��AsM
�<��� r?
'A�7s73�0�0� s's"���  zA<Us�H�����  �����1���@��h�t<�+t��z0���������v.�	��ӊ6OPR��A{�'�71�x��xv��v8lZX���  8.���v�*���n|� Q ����Q�Ⱥ � w�.{�Yp�PQ���t�  YX���s��[����X�XY��>
't��TV�;� �����@Y 	' nuSsX�r#�X�71
7*t�nr Ò�7�݋�  ��@<u�  ��ܔ�Rݱ<Lt��<{S}N�2�<F`t�Bu܈'� �^��
  �ZS[r��   ���#��U��t�R�P���03=t� �&�v�
& {���[���rtZ�5����-ހ� �H�� ����:���\���w?wK�6��»�vP�a��v	s�@1t���I2 ��&�t���x
�y�w.x.�~��>$��P3����G�D��1Gv ���FF���w���H�|ws�}�������P�+�Ɂ� wJ������ ���sSD��%}  �A�0�Ѹ�4� ��c.���' ����[D���F����&��X2��d����&= ������R78@�9t��uK�9Gt>�N�"D8Cju�u� ��#��6 �/W��C���C���<��C�B��\�Xd �.� %&�uX��ϰ  � X�P����!
��!�&�'
�u(�;=x���@���C�a!|
� ������Y�X�PL�
='��<fLEO>��f�����_��.CoC$�Cb ӎ�4���  ��d�" L���qu�\���y������x"� `˸ ��C� � '�阒�q��: �����z��D��}�"��\��r�p}P� ƍx���l�� �y��x=�$��V�%�03�Ƅ'x
'L'O ��Ǆ'�[��^�Ü�93��� �'�'�7�$`'�ȎغZ&/q�^� 4{%�� ��ȣ�&�'� 7'@�$Du�X����$� 6g���;R�>'�� �*����Ct��8�9Z����N�������{���t1J1��#�� n��Cs���u �<,r���"�VP,�� � *2����� ��Xt%�t�6�&�����""<�u�� z�c`�*^��&  ��> ��S�?��Ƙ.+���x~I���ܟ&D  �[��S�܋O[�Î �Ӌ��Q�Ϣ'��`:���D��r���'��<�;��!�	  �q���
�0�'��!�v� ��A:��.T /�S?p &�&`���]���s��LuZ�U=V=܋L<	�
t>�*K
JD�!<t:�
(靏�� �lU��r3۴Yz=  �=! �]�A�Q�v�T���tG< $�؜�&�'|
'>	
'A��ê	�|��L��|�q |����^4 F� ô�� PSR��BGx$x�6&'�oR(*	@,.'3Ҏ"'$k�����=��љ23�N�t&3��%�适��3S�f�6;�up
�&*

.�
�z*e[�����d�لI�
('�
,'p���Z Q���:  
��uW��,:�rN:�  rJ:�tF�%�>*�� D���Î��Ŋ�
 �j���ʇ��  ���r����g����
 �]��3iuUi����6���F�R6�\�� 2�P��ڣN�2X�bZ� >&����B��B:�v �������P�]7���� X�=�ȓ��;!�`M�+���Ru�>1�'$�SQPșR��9+�J_J�lP��U�Xy�0;it"��
����� u��'P> 	 غ���
�xZX�)�6���=\tw�� ��tn��!:	@u<g����V��| ~��6
�)&�p�"�]:tf rHEHˀ�ܝt ���	���t�����+�A�	����IGG�RP��.�� �Ɯ���ʋa3��G����<'�Z;hu��� n$&1g���Y8��Z����.̌�͂�m�K��0�I���-`:�t N@��(��.� �X���6��8 Cr��2���W
����t�I��t�Y@�����>����sH\�2� ����R�5���� 
�?X:`l,w:&v�\E 9�0'  Xu�����'&'&�f )�O8����03�r�@��:.TuL^����Er� qn>?�s]�97?`>?�Vv;Qk���"���W�f|3Ɇ�&��\I<�����M�����6��7�_6_-4'�>����2' �؆�:�u:�teS|�Yr?�t%��`�t2�:�u�Ę#� r.�:u��:Ou���8�*���>�k��!����m�d������QZ1`�-4��6.0�C�����	���'`n�Y�V��6F�H����v	�ɴ���� �$�� `��2�^��6 �:C�
�t<w1��
�$��w%_�
��t����l����
m�
R�K���� \��P6�6' נ:�'t��t6�O����h98'
6M��7Mt�2H��ē��t	���׀��r���7'����f ���� �9@u39Jtr�> DH�3�PR���ZX��4�>���rc��SRy GYZY:�<@:6:R����<F{ t��@ͨt�07BS�<!!K�XE@ ��<�����\������ֆ�:�p�9u�2����t.B��<`pt�s=�h��P�A觐�ڏ��#�<P�8�/ܝ� �K��)uQ ��U� ���Y���֋��! ���KZ��W�0 6<'SPG�:'��R�т23�P� �H�L'Z�N'X��3�0@P'�;�T'[�˻�RUsXǢ	�_��Q_ pS�P��6�'��F.���Ni+��B�J��Ās��B���b�
2�D�� �t#�+��0$�Z�`X(@Ȁ�?� �M  �ƅm�چ�MN:N_N 9
�  P�)T� )-���))�^ �n)S)3S'�)1)ꆕ�) c��
����	� �>t"\2�Q� �����(t�����)e�$�X�2
#u&� ��>�'@w<v�E��9S/:�(M8t�1�M` ����p�ñ��Pj:�t^qf���i�Y�t�HI@+t���32-�
��������� ���'��ǜ��.�>��g(�i�Wp�͑�-\ ���&�L���*�\{�v�(��@���_�|t�"@8+u��0%�k�t� �D!t�*2u�2�(�����1��C����X�Do��ã���QY�:' w
�
�u:T w<r�t�:��=. j���� ���t�<w����w������
#�ن��u �����
\��$���£ P������
׀����������
��	�&���Ȋڢt2����� �Ƹ  n�@Ո�	��M� ��ωP � !!� 3D��N�  N�N�NO���A�A�A�  A�A�D-EoE�A"BHB� �BO�B%C�CD~&gꕼrgי`g&�� g�� k f��z��g�Ag ;=? ?.��t N������g
�����$�$��� ���p=�$  7$fܰ?��\��(t
2�����G�t��ZG#�`�D%��;/�t*��� /�%�>'�=��u;n�tnS��� �[ZXr
�u��;�s��� #�Z3���������څJӁ8%Ћ�` �<'������.:�:'
6(8��6P:'vP������
� �;'X��D�P�@��%��<�u��RP�u�lx'�$�[�"�
3�

�)��������#a ��$������=�.���-� ��t���� B8�� c�q �
c:�v����
=`�(=��E�E�E  �E�E�E�EFXF�F�F  r��F�FG<GbG�G-H *�HI\LM|��g@�>�g\�Pg����g�g
�g�gr�SB�gMgǍ
�Dgg� ��_gI�<�g9G`G��wg-��g�zgGMg6G�q�g�	g?�g5�5�T5�g	�T5g?i'ξ�g4��g#�\xY��  ;=?�D������-e��	t\���|d�G��HG��8��6)�Ȣ,���/	t-�N./y�/�D/u/��1��, 3T�w.���k2��H>u�P�}+t"u��*A;�pI��u�+�#�p����ςj��Ps��X��&*ʴ�7��{����ņ�N�X���BD<l�Q	I� 3I -0  '�r��W����8�.T�_<��r
�
 j
PS��E�N].׏�.J��>\�Yt8"r3PQ�6:'yc�%��YX���tS3ۘ���r[r�>Q7�7q!�R*W	��� �����&�"�2�u'*��!�N��
�u�pOu�"�2����Z��E#AFzAFA�� ���sNx;6V'�no�;�:.T'H�  ����ݽ��2�Ja�r��I�0�tG��� ;>?؀u�&:u��u�rX�OE2+b���ah��N �3��Ǻ��2�VEt%M����"Ǟ&"Z?�a� 8���><'>W���>A�`�b���N���^_ `�t	2�����K���.x�[�������ʓz$�X`U�@t�Kt��s�Fx����ڋ��0�I��{R	0#�6B'V�D��� �3�>I+���t*�&M7կ�EG�&Ou�pZ,诹G�_WV�M�����y�r����x޸�\�4��{�F�yڰ �a��6o'���J��� ���6�>������ ������v&�%G Ċ�u��'���"�᪑���P��EM�6�E' �6"n'$�6�X�\e��O����U��%�$�R"���Y���Z�$Fn�����/�P7����P#�#70X�r�� ���;�s1o�1/w�P"��+�X�J����Č�����ˀ3 P��Äv�@a a����֖��n6�����Ǘ��$XG�&��H�g��ϻg�{�g�g��בg�	������g�g.��g�g'�##Q�ϗ�g�허 �����-�N�i �x���ј��
�F�0 ys�Z�� �	
D?D*�E*�O??L���.���:3^ 33$(-2K�80?d?�h/?/�gk���'/7D?7=['�=�f&?16:?��:61���1�3�����63m�l�7�L�����c�f���j{k��
�D=
[��f&����o\������
��0GtE7ķ>���P 	m���P����q% �%_����"û��u�_Pt�K<t��;q#�G<�KG<j$GDZ����B$�tDH�w���"n>|n� �9� �,�� h$3�3�D��?��t���P���1M*ۺa��� X?r�������Y[���w\c�ے��A����7����i��u�P�鐶��0p4��£<'Ɖ�H��pv��:�f�	�����&���F3 �sf �y� �E���6H'E��嫽  �Q!�!6J !�û�����  G�Ř2�����.��_����*����S�������;�wM��+ʇ�l����6nT(��)��Ft�֬wt��& �&���Ъ�o0G1\~�x�WČ������ [�3ҹ@��8�~���СP'�}VR�cKX'�R:�@!6?3�3��,tO8:� ¢�
�C��!1G5��SQ��Y[dZ�;U����>��5uKt
GG_v�O�P��->B'őBS_wKM^	^G_O��[6[Z)=�]��0<a��@���� ��\����   � �T�`�i��T�Z�4� ���1��
� �t&���Bc�d�$n�_Ħט
�� [*��d��H\��G-��d�h�y��
��% ���j�  �ܚ� m��$�@��a� �b *�����	��-!���@�� #@�t����#&�L	�Le#�e��&��ȉ�@}���w�t#\�r8�]r���mTd�"���#�3��� ����� ��؁>� �OLuXR IVuP �����=F�tD= �&t?&�&�U�Lu,< PAt$6"�" =VGy=E�=Gut;� �%�t�?�� �Ì�&���S�ʚ	�	���Qy���g��ᵿ*�c����8 �ˀ��^�xs%����
�x�Ga����	�� �Bx]� 3ɋ�G|8x��9  ��v�~�p&� �aw��S� ��R X�3�� �������s�w���}n������Dx�FG<y��w;v
;���u��W � �w��we�W�F�7� 0�P��v��p �VP�D�ؘ
 �>�.;r�`n  GG�.�9�ߓ�t'XP�ඤ�W
w!_��%^ �P���&Q� ���^sudYAtJp5�~�k��$(�m��ӿ�'��C� ��t�Q�YB  t���̨u&Bu
�}�`�/�	��Jt
�u��d(�B颌m��m ��~�N���Ds~�*����U�50��. ���V�n ���L�RP�V�6
Wv���=�(�)����^r�è��)^��)�� _�#m���$v�,�������jh�ȅ��+�9�V�v't  O�D�t����|��t����n��0�<�u<�t ��\+\�� <�t�P�K��=Ho�+C+2<��a ^�P��w���tb^��.���Óg�V8  u3��+k ������� �"`��d����0�� ¨���3�?uN�N��P�۴>�!X?�N�[i�'E� T�П˶��_���s��6\�����&o��Z�ހ&���^ �����f P��0����y@ �yV������5�k&$� �=���<&��K��u�"�~ � �`�X�W ��u���ǀ3<
��<Q��'lS�� 1��WQ� *�G$��PHr���: ����.�Q��
��00�YÃ� ��<9~�0��*1ux*��0*vL`�0�1����� ��p�����&�� �z'���C�>�v�u	  �$�{'&��x'Lx��%	J���0�����Lq��V�4
�t	���'! �2j2���33��3�IN�x�`9���t
&
�� &B&8K8���4'`$ɋv�~Z� *EaK��oNK�R�KK�2�K2�2d2���� �3�@�h��{o:�u�T��#����E�	`L ��@�R�D�!����V0��Mou�ic�0K��0 �Ei�X�.��.�@b�	���� �]iV�ot��������o[t��$�K� �u���ߍ| i�b=��VuDPQR�S��  )SWP����X_[��N   PW��f�Y����o  ��]���
S�/  [��ZYX&�}{^�V� @ �>p'�r'�
�e�P��;xw��u��h�h`�>�;������͉����`�� ������n������� � �� �W�O�?���O�DC L�
���L3�9O�31Q��D��5	��
 �w�VWo����	��Q	t����4�i� �r������u���G��x�L`�Z�� 6��#���x�q
�A,���)����3_�%  3Ҏڇ� ���' ���SV����~�t��
�'� �͹������� ���H�����5�!��D�`�%���!"��&�!3���VS�8P��'�< E��a`��G���O(����f0�WWX[� SR�դ��CC.���;�u�ZSK  �n �U�%,�X��  ` @ `	0 � �%#)K~0����=�Ŝ�J�� �l���D
� ?��3�����B� �DJ3�4	�#&��W ��QW ���3��>) ux��ԭ�6�u�|#t	�;so�DqĨ �E�s\��0sI` 
�tA��D�����îϋ��+ ���s�° ����u D��7 ��r��������  =�t���=2�_Y������P��1M��'0y�
�|  ���D�M����� 
�
��u� ������u���#	�V�!���WVRQ��w�z@z�P���X��t�.���'�;5��>6'Q Hd�3Ҋ����� Ǫ�[YZ^_�����R��XR�W�L+L{BzjQR��t�t�^�L
���Q3�����Y� ���Wt� �@#����G 0�� � �  J��t���&�'t�f!
��,)�"������2,�3ۇ�WNo�� o�WR.�<���Fs'���vQ)���B��X*1�֋���ܧ�Z��#�  � xX `Z_�~�S�����	'��$t���}� ��<t�E
��� �= f�w;wt&%�%O��

< u�E����E �0� 	�7�����&�-7I����Re<�"6�6��p"2 �D=E�}�D���t

ۉ o
#�@�U�l�Vt�7J�  �~� �:  �1��e���ਅ�8  �i�m�q|�y��L��V���^�����G�sX ��u�
�&� ��  ���_u����(t�
P�VXr�T@� n�pb�( s%��:��ڜ�s����<u{�ۃ� ���uEF.?%�3�
3w.� z+D�� D.�y0��3b��T&�@F�����\��!���P ���G#cx@^`R�
�4*bq�$���g��a�+�ЋV���$� �L�^쌿a�ag$�1� ֔ad����R��=�qɋ�S��1�B ��!r�[�`p`oN��RP��� ������X��Z�������
ÈTÊd����� ���oI��WiA�$�\;\u���&��\`r4x���3ۉ�@�D8�6�u���0N����.��& �_��+"3��8p���;#�F��`���`jg�CQá�V]�`;�t`H3tP@Xty@9�ZD%��`é"0�~t1S�JrQ#Y��ƞ�S��[8>�D�< ��T	ô@=��]?S�t�f�[]l��PQW��+��s�_Y�=��~�r8�� �x.u�*��<f�L�HxT�L;�@�P:p��X�DÌC��_T�ѝ'�E܅QP�XP�K�	ZrF� lD�	��u
�
C�^M x�) u��+�� �c�[���t�\̰%
Է����q�j����\1��4�4?�@��L� d���^�2�=��Ё���j ΋�PS��[r?;�Yr�A� � /�_I��3��@i�8�� ��L�1R�T��@E�\�@�Z��PР9r�Xå���-����g� ��d$��(���`��_��<F��A3�Os��| =hA;2�^�z^Id�(�= *�'R4 ��V�"< t�<t<�<t	י�Fp�L^�3��j�cg�s��=y{޺DDN^�NKۻ����` �д]�����@���:��<�Wg��W  �-@:��V�XR��賧� ��Z_R�O;�u�*.� ���p��. �I �# i��A �,)�>�y(���)�� 	A��|�Y�f"�PO�6
�� @��RP�T[����tV ;� 84t8 @t��-�����6]�f]
����r����bt�Sl��F2.,w��N� 8��H� ]�N�V��U�QRrK����0P���X^_�Ip&
�!-,)+���r#������YZ[F8�$�\ȚW0=�t���\�\ `>A��� ��&�W� 
��pSPX�+3�% �!�3ۀ>�&tFDCt�C���dr uX��uS�E�K�p=�9�4uXtP�%0^\=�u�����<�L��Fh�!sS(N~-^#�E�$tR�K��5a
�&au������Mt����[A��-�r =R
���[XZY��RQ7�������� Y�Lu�π�V���^[�\`p�� ���  �*$�D��� �%rl�u�D�y~��F���N�o�b�@<:�cȀ�t,�� �s��L������^���r��KB��n�6����X����$�#� �5
�&�ҋ<pô=��3��V#l�Yt��u��\�\��W8��u���Z�a_��^�}Q�&0 �t!�q�ك�R�0�,\Z����OD��fڀZ� �܀�����&��z
����.�r�^
B��@�O���|4�����o�Ƨ�S�_����`'��It@``Ot�Rt�NA��Bu�� HC[�BcW@�����W��wP�2��``���1�����P7�ظ  ��t'D�ʌ! 2��C�
�
 ƀu�@ ���D\9���s�)��.��^Z�Q8����6QZr$ZY�QX�   V�����  �_����;X"��~����~n0G�К�"�^�V����:#� d˯�������:�@>v���LI��I�^3-I�Y
p��cPR�4��#
Z��I�ޡ��:���  P�hw�X&=ˀo�X�XBی�0� �S��RV�J�< t< `=t���=+�t9It<=u���\��*;t�N@�_Q�9�� ��Wt,Q��t m+Y_���$X2 9�X��&��'+" �Ar�^�u�.���XY��6���cx4'r"��W;0t	n����I
�u���P�=l�X�G�,[�/�aaӄ謡]t)�W6��S��M ��HċɋҧrH5�`��g
d�m
� w4��V�Z�	UnQ��_R :�R��Y�u����WQ��x�@�����F
�+�I- P*K��`X�*6_0��SW�AWz sӞ��� w��W���J�]B��m�@�*Q�_Y�'��� �C�\t�����ͬi۹L��ꈋ�/�W_�4y� N��&˻��?(�u ��T������V�g9u�h���6�)�'�� !@��'�� /C�� ���|w;Q������ �h�_�� 3��Ǿ�)��=# 0���&8u쿾)BF����`V�.�P��3��8tFA�9�x�R�L�9=�:;� �_��	�#�E_�e@ �V�V�<�>����
����X"w� ���	#$���3�P�����C8 �.#���8��V��I��ҁ>�3�s������ 3.^ˀ&��L5�DV9�`Mg���x<������$���SS�����u��ʱKt���Û%�3��'2D�ҰÊ���8��e�ru���@
C������Ü�W@��R�w:�t�&	�A�R�f� ����M�F�����Z�}�X�$Z.-��B����K����'�iXY��3�v�Pl��'K�Â�'�! ��n
`$���@���'���ɞ�'Ro����� 0	��������)1����=�)<<  ��@Ɗ׊�����<@` u�����)׀��<v�PRQ���2 �0�v � ���BY��ZXP ��YX:u:�p�:. %����&��A�` ����u  �u	������p��ŉ�Y�7u��t�:&LRJ�᥀���0����0Ÿ�<r�*��AH�'����٥ 3@Nt
����7cr͇
9��fP���H�;��:4W���'�'	�'�&w��0 �۴��<u<� �]1�E-��'�=&����'&��'�{m�L5��N	� �rRI��8����� ���u:��'%0 <0D��:�u*()�(����	r
��H��.J��2��0�����:$0��9�	� ;wt�Ӻ<Ct�> w�   � "���RĀ��t -��tu @ M�
�.
�n%��_@8�&���n�uR�e`��&�&焀�0�_�$	�&�'��"�#�'  ;�N8(2�e_��d�W3i��Z��0���$,C��͋k&���u�3�0E����!K8���d����F	�	G&��'O&�'#�B$�B��.��3�o�kP��86�X<tw0�R��ʊ6 ;����+ ���QI���08�J�>-|���Z����[��A����X�~w<w�.� �8VP����9�}�Xe+�V�>���  �> t�3ÊEJ��q�JW�	 _B	B^��6 u5� bD ��6� t!R������\��'�����t������Z��
��0�s��	�B��Ou��{�Ǘ- ���&��P 6����� ��6 H�\'�6�%�NZ����*���2�o���u��.� 	����8�o�L ]R���r8�'t�)"�oR<q���0% �G
��-���V�w
�F;wu�Yx���w
&�
�?�OfV:"ҕ�������� � ���5 s�)�s��
��0z�
3��^ܑ���I� ���@���޴Hu.���!u��=�u�!�B�O`�L��'�?�%�0���۞�`Q<A�ģ&@: �\!I�#�J��á. J���Qr�`�/w���x ��Y�  (�������� #�����@ꂃ���� �! ��� �   ;!<"=#>$?%@&A  'B(C)D*�+�,�-�.�  /�0�1�AB0C.D E  F!G"H#IJ$K%L&M2  N1OPQRSTU  V/WX-YZ,��su  tGwO�RvM  KHPS�����I  �Q�r�x�y�z�{�|�}  �~�����������  ��)� P��)�r<w<  v<r
,��.��|�n��ƜUn��
&{'�Ep�u�t�UT�m �K�ν��C
�'�0W��L�� ��t<�t,<�t7 w�u0���2���<� Tr<rrn���t�:0`�u����*�r��pH��� ��[�0<�u�&܆�6�y`��	.ט$`����ss�t�S���<�{;s=��z��v�ut=�,	=���t	ʪ�(r
 ��u>����9%��%%u'��i$�. `�g��(�����:�t�-�����2�� �K ����:��k�b8tB����q���8��&�������.�;Q�=30Y�  ar<zw$�Ç���PRN�Zr�1�aP�<�����9G�N�)���Î� ~���J��s� �r١6@���@ ��ȉ )����� (ȣ�(9�(�(��)�)���pS�>*�
� n(#����j�L�&;�w�r	��&+w �r@^Ñ��0: ;�r;�wH�{�� �P�O���.�X W� ��Q�uD��(�a ��s>�t���u� ts0����+������,��>PS(�{[X�0}�^"�	z�zC����� �P�|�T�M M+���+�;�r`�G��\ Y��+�*������0���;!��v� ?+/;���3�|���S�^�������[�.���na�'Q�� ��c3D��_D_GO���]���v �������[;����lc%SQH�K�]��nË�+���{8��J{M�)�dp��]\V��r3_eǰ�9  ^�S9]WcBS���I|1՚��8��'�\���ڜ+ ��!�9Aw�>ރ| 5�	��_8k�MIV4s ���й N�1:�+�+ٷ@�ێ�r����$�3�0�i���u��4GGI���`#^Ì؀�Gl)w� �V���+6G ���A��� ;�3�d�#��lx�4�yL�
)�^�Q���u{�2 +�<"�v�SLs3���I0�% ��t���]TB���@(��;�h��W[��n���Tx; �tN�@ ����ޡr<;��d3��t�E+?�n������:�U <4�!2�Х��G�%+��V�V�W����t��X�@p6�[��]i�$��hX ΋��(���W�t�� �;�r�;�sb�_L��> ��\�	��;�u��d�^�nM�����6 �����	�L���'� �`) �|u�� �rA�y-�������v��@�8��Qk�w[���Ћ��!hh� �k+�� s <�r��+��h"[�5�"EɡGF��I��r]�	s;��:��=܄y�Ec��,v
3�v<�HP!O$.Ń�|	rF�;A;�r���"������0@�)á����S��2a�,���<��2���R�G�8 Z�< ?�ƴ�y  �d� � ��'�5��=i�RP��2]��X�	��t
·�:���Qy�Z$�SG�;�����U� ���l�
�d��ē�� Ĵv_�ٴ+�$�	[�aN���CL�
�4�MSR�*[��'C�-����� 
� ��P��d�r ���d�Ŋ������ӡ���D;������nfVz��frxC�2ҁ-b�|�j�u&u .��2r�ƀ�<`cr� ��l	��!	�[j]�:�`�oS
VwFG.y�{��I�</`�-u��:.u��������q�a���
��F��,  0r<
�rIF��
00 A�'C�C��ۯ��@M����V�
ҫC����C q��F�� �Mȷ�bu��h��%���~�����ۆ)�R 2�蓲�R�Zt�sk!� X���K��	) .1%�!��]Xô���&
r����z
P� � u�<t�R�끔U�
)P7><�u+4N<vC��tP� w����ƈ��Xu��S�Y� [��v=�� C�����.��D.du�y	��j�t�0Ɩ�/<5� ���<!s-q&Pp,<vv<  |<
SQ����P��3.�� ��^�� ��x�:�  ,�E�%��U�fʈʚ�ߎ$� b'Xs��fB��
t������ =
 t���<	r t"v���ø ����A���n�$�7@�#�>��:6�s��d0��v ����״P3Ҡ��9*u���u�����.�tॺ<nLu
-$!{�_�
"��28���s6c���˰���r�- S�7��  P�$�`�˃��u����-��u��w���&�&�0�C�	��!�9 r:
u�7>��ǰ��>��t�	ãr��:ir��t��J�J�����B��&.3��&ɀv����@�@�H=� w�@��:]�W���1�X�$r�����[�+S���p^�&2��h^���%2�

�:
��tQP� A����r�XY@�~3�� ���O2�����t  �t��GtH� �f�S:3ۊ���F�n�����)�A�	����� [��Y[�C��R�7�o�ՇW0&�)��ZYz�[R ?tF��� ��� ��$:� 2Ê�P��2������t�׻@z 5X�����s�@Z����u����H c��#�`�)�䰻� 6�? uQ�o`����u
��,`.I��YCJ��5�uM3��L���"��*Ș��Z$�$k�� ]�V�̰������ �S� 8£Kt.Ct3 !
Cu�6�w`e6�6a�+�V��u� ��>�˹�U�e @h����,�V�c�  ���ϧ��Єэ�Z�(��PW��E��E  _@������}���>����'�j �A'����;)���� w��A��tDC���nY�M��A�7~�X�U7��������Sb�?�ut@���E �O>�R>`�,�r*U� Ty� 3�.:�� ��tC���$>NOEMS�]�`Zs�(�m� (��r�w݈U�3��nwB�}��/"$�Ѐ 6�1��w���u�~ �r���=.5u����6O�<3�T��E�
��;������� 7�7��SRu�M��ɜw.�{r���==POb�0��1'�'�2`�Du�� �=DC�����=h�
+ �<�=B]��Tu	�� y�=FLuQ@�=I\�Bu{<Nu��;�u�ؤPAu�:W+e����hE<<Pu�!�W�.̘u��;�w;������P!!�M�\ ��<	t�<,��t���N��S� ���r'N��`���s ,0(w��x�<��ӫ W�s��t<[��á,#%8����N� ���i��0ދ�M+��$us��h�� nl��6<@d�B��<P
8����2�X��Q u3�c]�p�CK��4RP�����X��Z���-t�e�
Àt�d�D�	v4و�q�b���B�<1D��������!����b�
�[D��� \�%Q��Y�S�\�8��Q4�W�3 U_��u���	p�� ;���p��p'�W����� �_��/ _&�{�8��� &�9E�����#�	���/��G՜��� �Z���� �� �M_X<wF��g�/��G�_oX�5tR����u��ZG�7��i�� @� ��< r���:�r�qZ	�5�#���<	=I������0�	�<���2� ;@t�
��7��
u�t15�C<���u�Ms�m�P6�X�eÊd����& |��Ë��8���Ã� ]��)��v3�H:���!� <W��'�)�9��� ������h���T��_^�d73�MF�.߃ы/�<Hi��/ K�,o"
n���t24 �C������9͒5�P ��4��9~��=�f��XU���: WV�ꂺ3 9���ơ�^_  �u�t��R� ;U���Z���J; �L�l @���u�
9�I��8� =��U� ��K��s��Tp�*�b\��8�"E���� ��ۙ�X���Ҍ` E�u3W�xt
�tm ��L�gm� QW  �����ȾL�V�HpW x�_Y��_�"��~�s ��=�s��s�*虙��7���L�����"�Ju��
J`�9:�v�0�=vֵ:�3� �Iٜ��IOʜ�t
��Bڛ&��&u��ڗa��s�9�~� �� �%��) (�"��t螙�>n�y$�&n�  V�"�n2��0㘶�2������_�=	�� w/�� <��ř�e��7O��u��tF�p
�#蓙�v�.�cx�#��oc�c�2{,��r/mR��1�6N�  f�˸ P$�J�XPt����� ��X��<r�À���� NU�� u���Hd��$�r�i6wʹ$,C�ȗ���s��c�r�������ʊ���e�P� �� � ������)h��!<�蟘�:���!�bW���p���5\R�V '���t��	 ��A���Qs�d��r`�ZID� 2mm�Z��XZ �[RP�6� �7��:`��x��  �. 0��,P� ��� P�� ��� �L���=��p�����$�6�-1H3��g &�� ��-�-�G�M�7�>���t��
���m�q"�#�F�f8D@�F�P3�M�P @C^�An ���l 3���^� �.� X����t����g�x�w���p/����]� �- u�y'��T��>�-��3��;��=:-  �N� W��  �<&u[F� �<ht n�<otNS ��� Z_���s��@u0*t0 �	%u� �  "F���F�$ !�� ��] �
��F�� ���谞��_�-��c�� P�u��%u�$7���Aɀqt����1O#t !��%t�,���'p
�u��c��0���F�]t&�&t"�{!1�u ��9�5_��=� 8E�e��V��\���rr+�3��� ��U�<]
n�+Ҭ�"t� ����w&ҋ�  ј����W�>`` �	 �_�XN���^ ��� ��-�x��-%�<��-��-����@y-À���!������$�0 D0��t ,�}+��&\��`8� }{ |��$L�K O   & Q U \ Z s r �`  � � �I � � �   � � � � � � � �   � � � � � � � �   � � � � � � � �   � � � � � � � �   � � � �  "#;  @GHLb y e f ��t � ���  � ; < �&: RJ � �! " � � E�P�� Y [ J ^�  �C 9 7 8 � l n /�o:6z�N	l
�=hu
] I��T]$� � � 㝣�"����q��6D v X���7�8���Z�4&��# �  �  � � |� � �:t4�* 5ZfVL W�(Q*�@$T*j8�~fQf�^�Nx*:t�Z,��2`hMY48DL��>k*��~�d XQh��zQR�< �T�(�E���~|S�V=ZX�"�m� b

�*E6h 	 g ( * + ,� m fw�
��%(0*h~� i�(p�@8>` �٠$=&���� �݋:OtF��� Q�A�. U�����-�_
���=�5�Y�I H���7�Ў��")M-FF,�?��.-  �O�X+G|;G }���ٓAE���!�	��D��D��D�D�JD�D�Di�!?�7�$��!�i�F��]cg�!h=�V:�� V~�=VV�( VwY� ��m���S m��mzrm�m�5�h�> ��R8�$�"=��ABxBk�B��Gm��~
m��m��u%mm����k�=�dh,8o�$md��AE�EA2@m9E�_��F������=������k،��
��|،��]��iS�)t@�
�?@�)����ՠ�c�-�' y�RS&�\���Oq����U�������
�Ԅk�k� -k~�l��`w�l�
zjl��E?l�,s0z5l���5�
�ԃ�!/'tl���i�kR���Y���$xv���C�żS�*AS4;��6D?	���-������5xqq��al}��=� � J�3��G ft@P�O+<f&<<<<��<3��-/��f-% ���r+� P �R���6�� Yv?��*%  t
<r	P� ��A�P�� P�>* puYXQ�Q�@= ' L΀R�6
�xp#���X��� �� �Z �XR�Wu��@t�<�4'9t9��2@� �S����*��V�� ���B���*� �{$�<t�pQh�0 ���%zOu��K*(��yP=)�*iW�	X*�  S= w�).� [�QRP��TFZY�3��I��i���0�u���-Ё�
��ꢈo�m �O	@YÃ�8t�0���_�=m@"������t@IuB9��5���03� |%��txf������,��W����"���Y_^EY ��V���W�}���P��u� �%�ыȭ+E|���;}��JXHy��g NN_�Y�/���`���5�AXZRP� �
PP&�4���� Y���9�,
�X�XFF� �
֚Uc���R R=:G:�������=	��+qX,��-#I*P'�����v	��ucI�X�\�&�q�� =u �r�>j�q�q��az,>��c�6IO�t���0����B&N>��3t\��1=2��e�=�U���N=�v��$}.������
�0t��"���Κ12���.t�!��q�oл��Pp�PG��j
�܃��*,_3ۉ����u����6� � ��AW0fO�,:;.�r4^]��+�x v)W���)�� ����+Β�6�+�? �Z+���� �׋+�v� ��+?;���� h�w	�#�� ����@�\��-�I'p� s��#���.��'[>��&
����.��F����X�9z���}�V���E� A뤰Ft9N��ZB�9)�UPX83Ɇ��&�ra ◡E�968tn�	�x ��M��4p u�7�X�<`��C `��О!AI=q ���@�� �t¸���F�|6�F���A1~��(A�P�t�/�P�m��m�)��w0����l�\ 	���-&� ��c�-*�0`��s m�-����2	ݖ�;�_�����o��%��[��2�&��=
�+���OO� p�À�r�I�˳�?�z��w!($X�̀C;�w�PQ��d�&�?�#&t����%�=	��� X�D��# ���;�=XD���YP;ʇv����&T7&�~{(
tI;߭jb	'�z����������� �9�G�7�{��>  #�% ��X����$"�k����5]�S�9�% {b$CS�F$��� �9Z� +��|��Xi��q�܂�'��()�c!"-{�.��/	�0�1���28	2���#z  ��������9!$  '*-�6"%(+.�7 �#&) ,/�8(�[�-P���+   ��[��t�P�\#��.����[8�#*��&�,��\ s�	�3� �W#�##C#�D�^5^��"�� �"Q�"R[XZ �!#;
��"�J�@B��E�tnu��ECF�$�RP�"]6��"\�P�n�"�=>�"N��i�Y�X[@��:�� �GZ[��*G��@P= �2�~YZ�<�$���"�5_���4[鸧!99_w�=9 f�[�@p�;�V@FF�; ��%9}����,��[p��x�t�0� "�[�p؉�RQ���w��8���G[��w=�5�h�r8�0<Xf��4�\5��R>:�=�7Ky2�����E���S@T ��voG9G8=G9G9G�G��\*F������7UL��[�?  &4��h ���i 3G �
�uK��;0 �v�'0��u��� (���P�=�����Z��X ������-CYp�V���k�& �;&� v���o 9	u�^Nd���R ��ST6�������p/�/ gQ^�Huу~  B��-;FtXX���c�� jq�q>�<��w ���d
R�X�P0���l�%��j��-��. �B�Sx�7����+��-q4�'�3��R��q��II+�r;6�w�����.j!PT�2 �P� >Xa' Pb��?���@��L�~�� ~�� �z�`0|��v|��'p�,\�
{�H��B�4}��� �� E��� ~A�� �
=� ����� ��
�p���<=��|� t�1���S�>���A���[��S��>
p �y�4�a蘍�`�d�.�\.t���Aiem�i_��n��R��b0v��D��>��8��20�� =�	)��#N����yk=�x��D�������.��._�(��Fp@n�1�
�<
=q���8��f9�r\�A�TP��7�G@(顽�U)�>�c��9i��q���KViS�a@a4jY,�OYQ�K7	��#=S@��l��jh�G�hf�#�fd�R�P�t���Ln�
���
=����sRє)r"99bO���]��H�`1��{9Y�S���g!R����u�����'�S���Ilfo�}��B�A�@]��P����i�op��4	\���P�y��@�o?�����;�q�s%k�s�uuF�1c�
#w3���
yh}�zx@
�;�VP�%�
��YV��
��'�
��}��p
�@S�X��41��2
#��5�w�� ��,��+�f
�'S�	=����k>�ޟ?�y�X���@ps=��@Y��@CSK��I6:��O�V	����   �s}af�	 z(cHf.M]a�{�A�y�t�1�&�u"�t�" a Y����3�Gd`^"��.�_ 3�X����{����ght��Z���@Z4���'6�I�K ��=F0!PL �,y3IbJIb�$��P�ʍ 9u�����`�� �b'0�=1�q<�BMA�OG�`���SPp��R W!����	��9x1wP"�`3#k@.0`C/ZDIT�T�%��  �o��P�P�c �[�_�S�B�<�ą6A�0>�A*ʸ`�D!f�h�B
p�		I��Vz��  ����u����	��\����]�=+tC~�^���_�"������&4���a0���"��� ���Du�T PV'@$���vc�`) =� X�	��Dd�R�O�@�D5.� Y���� 3�Yj0o	[YZv���8WRQ��n�<p)�t��˰��t*E� �oɢ�ʐ#����]�������� �`���S��w 2��8�x_�W�� ��$��0���[}z�@��� ���\	�rd�U��d���~	��"�<��r ��"��d���d���d���d���d!���d%���d)����r=d|�/a�W�2�
%Y:���Sή��R����Qv��P���O���N���``M�	��L�
��g&tKie����s��k��<��x��l���f�h*jf-�3�0R�emVP� dk X� ��p�w) `�pYX��p�e|Uf`���3�l[x*�@jp��^o��_QX4�SkQ��`a���3�+�p�3E'= =; 0Y3�;�uKS�B��qt @ӏ,a"N�AKj|�S�?_~8+�>ED}�t���q`#���"u�	�y
1
�~����� �a��p,y&=�qK  �[�t_x@�ZH�W@Z�A��P)w)��@*p��;X"r�>�/Bd���u#bE�y�u�� p�4�*��I�V��x%!H���i!!H� �u�	���y�1���ZY[��3�B�a@������XP��P 5���rD�1 w���w'�6 q���s,�0Tk�� � 0���t�  �0Q��A ��@ ���:��8w��0p���(�� sv.�qɸ(���M�,����T�.����O1��̌�0&��$1��!�x������K���u�KrtHH�|������um�('U���#:f�M��w��
�A)�s� BG���6w6� �e�$r�s$� n�Ï>������	�gc9�&Z���Tf�eu��o]�\H��BT�Sc���HvK�J���t?���>B�u6�5ސ�9-�,����9$�#~�9�7���9���I6	���qވ <���`8��r��7�- %�0<�3���;�|;�*^�*��Z
��rLP
�����+�� �0��XwOCr~��� �X��uû�] ��$��OS��G" ����-�����/;w�s�Mfu�� -�G? ;�t ��&� ���*�(�(*�B�Rː&��X���R���ZUD���-�=@xjq�6� ��%3����k3[��	ǆۧ�Ne,T���؋N���� fuQ�B \= XTffPLHD�`@�>'n@阙-� <840��,($ 8!?��+� ���uCC����.��#�$ !���#�����$��@���6�u��@u��M��"r�7����������w��� �k���b�& =E����j������[�1���X�DM@dG���P8$�U' S��t����$m��m� p�� ��>�d"]4��L���5����
ff !"�Df.���p9@%�����|��X=ff����&���#v =�n�� 0�H3B8U<Y6:0;�L*UVޞ 0�(�"���իǮ �@s=�	?� vh�P�lk ��SP u&�:�)���к�g���x��~7!� ���A�%{�:��� �<��k��e���#��0�x����L���FxP��@��B�x��e��B��U���aA���R��&"��)�A�t���X���`��&�6���*�<���@�^���F�����?�Al�똓 #^t簖� %p��V�� )X� �r������� _�K���Ê��NҎUF�L��h9 =87����@t�G t��� X�X"|���E�:tF�*zV ��OII����+�r.;>~(����
3�  ����w��̀��>��g ��4��F�Ș�&W�"� �S�+[=G�[�8^>����>��E���+��5�r.DG�% fu	�_�h ��0��@u"�O����sv3�W	�EN���t1�	7
p/��
���U��I� �9rt@���8u�&�F�Ð��������w��+7[�2bS�2���#�
�X =v ���8�E��x�-�&�L�����II` �G$<m��<r��to9�t 0���W�
�=OP�Q<k�F �q>	2��� R@ŗK�gP�v�	tɌ�N� �2��X��^��v���n ����t'�� ��	�7m��
��w� ��t&<t(���  ���GG����	�i�NNKVUh0�����D�뀠DD��֌�V6�% �?�� �
 �$��,���
�� �q?��P�#����D��
��	œ�g	 �S��P��Z6ы=����� ��[���)�H�v�(
> [PSP������, �&l
"
9D�g�4 i�y��W��[�$�+  ���Ú�R��   c@��^���=��-[،�0����F���M�+�_^E9���P8ɆnX#����*2���1��M������W99w��Z_0 �_�O��Np^��?���/��Jiu������7����ko�}�7�����x3	���k�� �n�[B��  f��S���X�����+ l���s��6+�f`�ߎ^S��8 *���-�V��7 r
���ת�� ���{�}ܭ�бӆ����;O���L�K���Í�?��YPQP�qϜX�����B�+�ډ!4�%d�� �sW�'�c;	sKRR�	�N�X[�_��ۀ?�<��$��=�0��_��Z[a� QSR�F���?�X��ZXPߑ&�ݒ����3qnZ�Pw�?pQ7�4�^r��h��1���� :��>�oY>5�{.W���P�x� ��� '�D��p���Xk�HŭLȃ�F��v ���M�0̨� �=��!��3��������� �j�a �k �  0 �8���	;�v&�=���Gz��0�:�G<����W�  w:Ft
Nw<���R˸���N%���!=
�u����5_:b\W��Bu����^W9�^���m�)e�]"�X[�SQ`sPQ�K��Z�PRP� 0��,5!6@2u�
7	��4 ���v6�H�R7�I8%'�I�J4� 0h��G9�%J�K5����Ep�0	�2[��%S=�<$�`�d%�e*�zjZt�l-B���3���-�`B+�t2KP�=3MF:M�`�?LB9�E03�F-�N'x�Q�h��Q��Qv���S&����Y��C0Z�Z� �� Y_�u�L���Đ�=�Ĥs�_[X���ZSWPQR���T
�Y��� ��� � e�6������[  "�z6|A�7��~# `b JE�8e8���" @���%��$m ���������  z�}Ԁ�������n�q�  t�ec�8�G�&ggg  #g���f��8���%  ĭ�;|%Uc���g"d� `g>gO�g�8=Ԧ  s�7ҡ��/8����  �h,�h���%"�?�U�~ 4��(J)P��:�c�c  �7�j0�$�d�e�ct<  �?t��6R�Rc-e$R  tgqg��`8�,K,-d, -��Ҍӑ�.��Ȉ  �^�*��YR�`�|�@[O [:0R0^[�ZJ[Y[  �\J0b0h[�Z�Z�09?  k,01Z�Zy?*?E[T[  B0Z0c[�>N�w���ˡ  �a�a{#��bbb�� 0dj8&a.a�;�a�I  e�,H,-a,Fc~���  7�f>��G�ļ��T�  vxd�sũ���fpee  ����f�f�d�d�g�g�  gf���$�d�^�dw.�  -�.�Z��r/�.]�k�0�ҵo8���k�M$�&c�
� �a�a1�"?���f���f�8�̺�8���>�� 01>�=�=�=�=G>��>]���{s��  `=~;�;�;B;�=�9� .�ӹG8��A�M�N8 [.�@�]�O�	�U�L���WJzXZS<<��N �	� `��F�JX"�u"�4!��.,�,�&VC���}�! ��.���5�HQK��.
�!��s�u� )�-�Î�-� �,��e��8.ט�+  ܋G
=�,u����g���;�u Bm=�8s`��� ��0�!<� s� �=� +���0  r���ׁ�ns�0 s3�6�
 �:�}��0�6�&�� 6{�H6� �R9���+��۴JP6�} �f�, ���=� �� c��:*�ps+�Q� �T�:�� � �;���9X")3���! �P���B+�=�� � 5�kzm %��; 9 �"�.\1�}�6� ���"��3�6��"s)柟6�}�Z��/Lt�x7�;;�6��3�&`�v t,���^ �t����u� �o��� �����7����̃� �����D�r
�t�� �@Ky美"�� �	#�p@�v�.�VW
���,',�H�|'$'s �feR�	\ ���:����~��F�#��R\t�_^�e	s�L� �� ��k��H%�>�0!�� D � ��;�s�� ��Et����� �����<����  V� �;�t@�t�3 x�������떙���~��ƭ]�s Y� �+�r;r��RQf�ˡ@�7ul�.w�5���: 30ne�
�v��nË�s��m�M��3��c߃�u��A���$x��(��u���`r�s������bWVS3��b�}���ff74��SU
7
u�N7
93�����PF9��>��V����o���؎u��`�+RP�v
��\;%wr;��)v�����t<�ں� [^_��:�SW�W�������:cuG�L�)��f�+F
V�JG�_[�d����	6��n2A��� �����){�  M˄=�  �WU�]�_�E��DE �yD�D��=����=�� a$��.����tE˙X��\�� ������;^��=X��"^�zZ�~� f�t
F;")�H$��`��&���[VW-M︳�ت�{d�5�{lEdDf�����؟w��$�J ����b���z�a&�����������|� ���/�$ $>!�eP��#X.  ��>��6�Ή����3�  �A��
 � ��?3�$YY��� 
�+��u�� �Bt��0���.}�$ZiÉ >A�t�?g�v�7$�����X4�&�	X�u�ۣ��  ���t�ǀu
>��\ �6p9M]��� Ջ��r����3���6��������P�ڀ� ����� t��� 9�������X u[̀�2�3��� �toN<Dt@<Et3�> ��t_<+t<-uWN�$<� F�N'�t<9w<0r ��X�3����������������10/������n��
Du�@6`��t���~ܓ2���>

u l+>���:~��	��}	��xN�>�vN��5��7dt.� �}� Au"�>r�`hQ@y�mYÚ�9�A��`;���_U��K�ߋ׋��zr9;0	������k�D X�Z��� 0 ����r��Qs�X ���>@�xH�4 ����{\XV p
���������^�� WUS��� � NX3 ���������ю��#@�,��)2�3�A�)
�y )� r��)}�P���&����
�[�!!&�r�X(st ��	2��� �r����w����`p�x���|v t	t$$N�� �N�b�,0r�< N	~,r�
:08_}�20FN3��&%��(u�l�4����G%u��$>�x�<.t�B�Bwδ� �˴ �
��I;6�sp#��>�< t �,4<
t�<t�< �ar<zw$_�2��f��r�?�� �?�2�0���@�  ���t 0���t
�C��I��O� )��؎  ���&W� �^�L��d>�D�Kt��y�-^l���N%S�W:��Y��9 �7<3��-����  �ȺM�⑰M����x ����������C0 W�߾~���B_�D<�/�4U�VA�G�R��B:�W\E jy�����������J�?�ً���s ���������  �֚��ٿ3�� 2��UVP8:���֟��^�Y��Y����] 0��O I�0������l�Z[nz����  ��= s4��t `0�����ؙ����� �n�R ��/��v�����7�%���_J�H�AWI5�	 O�Gs�=�7r6 'N�W���Y���g�_j��a�pE����[3�
�t�y������������ 
��3�A"�
�� �������7딸s����R�	��F�
��5n����� ���� ��<t�� �^�<u
��u�lO<u�s�<	�oVks���@T)
�
�Q�
@�
P�D
$�
���9D
 ��
` ���4
������  N@��p+��ŝi@�%�  �O�@וC�)��@  �D�����@զ��I x3@����G���Ak  U'9��p�|B������~ ЪQCv���)/��&D�
ףp=  �?;�O��n��?,e  �X���?#�GG�ŧ�  ?�il��7��?�Bz��  ����?��a�w̫�?[ �Mľ����?S;u^  ���?��9E��ϔ?��  ��;1a�z?Y�~�S|�  _?/�����D?��9�  '��*?��d|F��U>  �#Tw����=:zc%C  1��<�8�G�� ��;�{ �E�y�9F��W_��F � �'����`W% t�S����
�2�� �[����5~��^����8��^�
���}R�V��%��F�  )N���������$ ט����H�����'B5�C�hn��P����Ŋ�P�&�]��
�;�c�?B6��5 ��RH�Tʹ��
� (#:���F�uX��7.h�~�a�
��X��Bt��
�uA7�W2s��
��� RN.�to���@u2�)19�n��;>�ܡ� f�-�?rO=@ sJ�w�����" ���I��� ؊�/"�"��tK
�V���`��5��y��>|�/r
�'���T���5�'Ҏ���7�x�R=�Au��#��\x����������C�����Xvp=u�� ����u���m��������j����I���R��uD�\�V���4�65�Ñw2������2"��P1�4��:�
5��8���/�����'����(ZyF{&X����[�{�_�&B<�&tŵ8J�?���f����.:�>9�5�'��1�����!��H� �D��,		�D��Y C*�; �R��H��������4р������
�t�r�QM��t��(
lÕ;����M�c7�����X�2,���Q�K#R$'�����"P���&��{�� tP������.��x}f�1`<�u�R ��+���t�E��I⺱��S2@b��EB70�)Ǩ�v3r[}v$h37�j��J�^髁����D�҃�
u�I/7��JC�����>�FL��~u�EG�F�p2	��l(E���#EL�������or�ƪ-�.>�fm@ʽ��Ĵ jWV.da�3۬����Pel�<+���9wa2�ҋ�H#��#F'��X-�ued4^_�QT�y "~
W���
�tF �
�-��۽x,\ÍU������0ov '���u�O�� ��D��D;�r�Xz�  ������ l�@O������6@ B��PLOO �RPDF T� 
 ���BB �3� *���RB����R__�@PEv�B@@9 @�t k߀rO Or�d8ī�1�T�[(B8??��O3�=h � 7����vE�� l��� 	��""�/	 q04b��Ā  � ��-@� �q6;�-nt��6T@�ÜS�J-6��At���G[�  *�&�D�P/�&���D��u� ܸ�p&\�G��ܘڨt�  &�8� ��� � ��p1�&��O���j�EUEOEu�SE�׈ �WQ  >&��n!&�|tb�0�[�G�t*�� �L�>�EQR� � PP�u8ZY7�T��(�&��NE8G�b��Lu���r ���� :Ou�Iu�"���u�H`�u����t� �
���O���� `�v3�r�>� 0�� &����i�
M�j���`?0���Q�`f��.��&ûj  � pQ�Y	1
  �r�	�	]�   Y�/	
3V= ��H	 
L8��6�
6c�4�
4X>2�
20F�
j�,| mN�V	. 
o�	�	�ZV�,	
0 @� E	
I�mgjd6�
��0 ��4�
�����2�
MPSJ< 0�z�,�,�,�,�x,���/��  �	�
���1��  	F
�U�v	j  
�!,n��	�
����>:|���	�
~��.�� �	C
�R�sx 	g
�)k��	  �
�������  &�G�����_��� � ��.��w�&��  ��&���[[������ ~�ɘy�.�=
�W��P��-��w��Ys��:�v��/�5[&�\tՑ�1#Z0 �)�)  �)�)�)�)�)�)T)Q)  N)K)H)E)B)?)3)-)  *)')$)!)))0)�F���P�2
�� �׋�GG����=�t���H��h��`����$�O���` ��?OO�G�>`R-���2��6��z 0�-���u��Fa8��5j ��&�D�%œ �" ��E� ��@��?uRP0"��3��ZI� u��[�&Y��܁X� \tbʀ�&&���W�| ����@tV�6� ���4^3���f qP��?��p;l r��0t{�R��� /�r
��������ZX����<X�vCrx�m7yAR`���-�F�����US��~
 ՍFPS��wE[  �  ZY��]Q�H�Y�@PQt���CC�GR�y��" � �E��p�	 �_t���� �D�2.0�7�,'3J��5�ž���N�P�OF�tFF� �z3䌑�<Yu��q Y�ޭ��� ��I��/`c���r1�	 ����ӊ� ��y�u��A����&��&��- sr3�=@3u F�O� ��-��0�p��p�a-t-�#�$+}+��N��Ka+J#uX4L8R-��Q&f �
=��sS�-� [�Y���b C��;�u>����Ӌ���K�����t#`���;Gu���=8=u#���@ ����6h4�%�83t� �� NN�62}�ð:HH'���r��V�� ;ه>� t�;�u�3����R��4.�Ǝ�1�p;.ֺ�S���
}��l�9Ls�E 귀��;�w&�=&���W&91�uO ���9>�t���wZ�� � X%�\�*@<rH pP�)XYW&�&�}���QQP��2�M̡������ݱ@�		�� ܁?R�Gp+���� ��)��)QS�رY�= $ ��� ��%1�	��2Nɋ:����=�������_�f��
�9�t' ����-HHS��6�� �uY[�t	S��ʐX�0[?u�0 |�DI*���r3�G@@_�a�K�[ǃ�I��9�lK��� �w
����pB)r$���?���y88�1J�����@ B0�H� ~h�OE>�ldZv��0���'(�'�.(H$
&��'E$�&��'Z$&� �'�$�%<'�'l$��%*'�'�$�%' {'~$�%'r'�x(��� '�pī��	� ��/  ���P�5S@t=HBP�UPP�   �� KK�7�����&SU�Sh�S�^Q0��~�Qs/2�p��E��:�sD�
�����u�"��F/���� a%�z�A���������p��u!�����Pu�$��#3נk�L��X�m��,��3^'��> u���W�t���!����$,�u@��$B���Hb7��'�+uI2�5\q6��ʫ.u���?%���|.���V����1o����F���Ê����&E��|Ե@b8�. �r@;^ s�^:so�:�t
�? _u\�CC ƃ�w!;uL�	r	��?;Q>	+�D5�^���9(���� t&��-PSQR�A[e{1�˒�N	P�����-�µA�w9�~@@�HH���1Y;�Yunژ�� �}+���� ��������2��  ����_^�&�+��M��: S��Xr&�a U�YP��ar�W'`6��F��� �'Z���� �)��_��+k+��@u
�O���w���t
����#�i����X(|�N2W�7 2G����S
u����@$�� r�3��A��f���A�=/�+�t��Դ��%Vdt�t	��TP��� 0�m%���O  ,��� �*�*�*�*�*�*� ��+�t-�s*�  (QR 0kPSP��Y[��@�W��q��_[^�ø� �	 ������+���
��Gk�R��Zu�8�@t�%���� }r���r����$dRQSnr��US�Kv��[YZ��kNNX�P�j�&�\��B�FF��s+��xuP�f�%�e$4�t��Pt�O:��O� V���9�DF4#ɍ�� �5 �sqT}\~T���W��������r�_�٘���봫%�\ ��E��TU��E�� �u	�g����g��$�&P�6�G�����މX�$����S �WS��s[�� PM��GGF�� �����0<�u����¨gYl" �% ���;6�̌s!�C���� 3����lë���	\���	 ~� � B�XYS�;�[*��5���r�����% �� PSR���& ��ÅL�M7[�J% �CX�� :�u��� t��
�:z:�t�X>[�B Q� P��)&������^��d�� ��� ��a��7>��l��lt�;��/5�
� ]�Ҙ�!2�����X[P���k`�v��H��
��ra����RW�� Q%,���i��m��c0r	��p��	q�  ��È�����0�����	�Ӏ�] �Q��(t`l#�^&+tIN��� X�( �Y���C����]�F���P�&�h��<O�%P�'�!�r��܋V�1
J���F%B
I?|.�}8u�G�N%@tH &:Tu�/��&2�l���$��PS�� a\O���	��-;���U�� [X�eG@����@@[
�T$�]"��:\�߃�=_�>��  l��3�.���5�j�u���� ��T��1H�'����P� �
Nϸ���X���<��2;�R�)��9�5�t��?��u�͠p�l_`  ��3���Riy�  �z�����#  T/Cr��������UQ.=#gU�$VO(e  ��,�\ fv��w� 7����r,@f� o������` ���6: ��4�$ilc`2L�����0b>�,�,�,�,�,h9�.��97�D� @�@u���%� !��*�������T&���� �&�\���u[S2�8�bqi�`q�  \q �R��Q��Z�3x���+��_H�s	q \%&�X[S
��  �����6T r��7J`  v��!���� ����������3Qo�9 �X4G]s�� �������� ��Ѩy�u�ׁ��7O  	XY���PWR�������܃�����`�k-�`[Hu
��s��#����2r�8�E��� <9�3�SZ� �P�;  �PG�uR�A�J5�oC��C����@:�� �Q$��t�z���2����P��s�'U���jL�t�=0�[t#��WY����X�����
k��0��W�D��#�'"�X/�1[[�B�1 I�H<r�ސ3��V����m�������j� � �� g 5#=#G#M#S P#Y#_#e#k#q#w#����
�6�=�%�W.� ��%�)�P���2��x5�а�xB�4�P����(��u�����X��� 
�S����s!�8��[�_��b���K��O�G ���	�G2�y?Z�Ku���L @ x#��u'q%p'7:�`[ �G��� �� @��"���eN	֓6��^�����S���-=�w	�<.�� m�6���It6;8V6�^��p\&GC�) � K�XPs��p�ܸ;5�	x�H55Ǽ��WPb�XZ�Ȩ�̫Wp[��@��g��E��Q�I/���j�\�߉�� 1B���]� Ĭ ���ȟ���0 �Ϙ�;�8�	y�A��I�x"�#���H~@�������W�mQ	1��t��۽��=�������2 d������ $����P`�L���cZ�e�h4@ ��S2仄k
  �x�2��	555%d5�*���*�"
�"0 
6�+�+�+�+�+�  +�+�+�+�+�+*,0,;��,P,�(��f<k�������� ��#40 �4�4�4RZbj��a��i^r�Xx� [�)�)�)�)�)  *u)�)25�m l�?sF(n(  �*�*�*�0�*�*N   00�*�*�*�  )(/?.`�f���  lru{���z  *�*%/�,�,�,�
�
��
�
���
  �
�
�*4.5 D< I F , ; -^x.8   {.�
����( �.}l% 
C TL��_  4:3@3� � � �  �"�lm
�+.�  "�"@ 48��":*  &,� ! �!�!�!�" / �c,n,�+�+V,��  �*�"�*�2� � �   +JQ�E!� c  �*+
33l+�2 $+N!T!Z!h!ry�.)
!!+��  ���"!"!A"y,^)  f)j)`+f+a"h"q"x" ����"���� ��23v  !|!�!�!$3*3F)�*~  "l+b)(!�"1+T+r+�  2n)�+KED" 1!9m�?!�"/  )4,�,�<�<=�<  �<=�4r&H�4�*d&  b 4*4�34
4$4�*  �� �y&�  .=�� Bh � � �   �4�4&=n �4�  4�4�4� � �&t �4�  4S4z40464<4j4FC `z ���2� �  � �4�4� � � L  �< +Y&5�&� ��   �k&�*+&A5G5  <xr�<�<=�<�< �<�#�#}#�#�#�  #�#�#�#�*=�<�<2 �#�#�<�<�<=�<�<����+�*V����?���x [��	���'��'v;o�aK  
&"+R"5"s0�|\6� Y#�;���&�4 �"�#$�#W	h	_� � �"�����6`8r#�C#�	0b&#`�"D
������F ~�7�88��
�&	�@�"���|ɚ�'e
�M+ y� � ���\�2���xy�
"�	��)|�j)��*�!+:���*Ea�X��s4�.�L�XXO+�@x"��&*
`����P��H� <���[���t��#($�J"���+���H(�~`�J+�Q"���*�^��9+�+��NNa� �F���o&�9�� !/�/�/�/�/Aְ%�P_ﳠXRӺ5����-NN��D��M��ap!ғ0�u �?+a� X .�[�W;�����SCFF���������&2�m�� W� ��XVW��  �2��N����&3E�%  �uY����% uTAtCI`�t@�����uOV=E�a  �C��w>RPS���,��sӂ�I��I���΄���|��Uv�_^-I15���+�B�� v�+����P���X߸yXY2wa ��HH+�;Gu�G�g	� �II�O��	+�ͫ�X��0�����& �t���pu�t��&�D�";��p7N!1�r�>0&70"���PT-�/�2I"d�D��P�xX@���2W"8\�B��V��-�OǇ�	�tSrP��������10�!�XP��I�-/W� T�Y�����"��P2��9�����H�2e��0��%  �����>qu�%q��$��h��ю&1&���]�Y����n��� a�@@�O���_-��'q�_�FF�7�6�^������T P��!�?Q�X��2�տ�w���@� D̊�% �=���u	X�.��m�1�P��0 -������o�	  �ً�&����Q��Y���h��ޢ �$�P��݀��lX� �u�C;�-u����"���� nr�"�3^!�
	2#�G�&SG&x�ZP=� u�H�e!�^�5d� ���K�:W�z� 3qX�W��S�F�0��&�5����(n�&t'�- 8P�
�y�a�@	6�"��5�@t	x����X�EV8�PR�" �VBu���&�5���J��P�x��XD@N�Z�� u � �"��(u��0��#���)����p����Ǚ����G�O�A�ĀnyH;�t  +% �΀X�<��������@@�Xh[5�T�0�2���&�EQ�� ��5�> �O|P��XY�ċ�;cX�`�wX[ϑ���� [t
P�-/�$U���L" ><��6I�t(�R��̽S�j X5Pb�qZ�N ��Q[�?��[���? ��Z�2��IK�*6�" WbW�$�Pz \u<~
<@�s�U��4  �&�G�-+�BB&�WV�ø"� �&�;�t*�Ӌ_����k�ܒ�����u��y!B����  ;�r���_�S����2��ƀuP�����g:�|��
��\�!�t3YQl�B]�@�[1A<�Hq��R�)�f7*:"�t YX.�tnfu)tiw1&��g]�uN '���&J�P�%uF��87��A ��D�X Ã�s�HH��/ ���tAu�w/����D<��j��?Pw�Rw�r� � RQ�fYZ<��I�$| � 8�X<u
��/S"Jp [�����g1�놋w��N�|����G�@;u�� ��)6�g�w�;�t#� 4�y�� ��_��F
��p���L�-�T�����َ�ÏF�L<*(1�5 �����X�� 
�-���X��e.`q�.���R�l�ڑ�C A��00)0D0]�|0  81l�%1l0&0A0Z�51|0v0y0s x"1�0�0�0�0�xL1�0�0�0�pI1X�9�*� ��= �@v�PS��Q��g�:������̠���*�>'q�a%���
$qu&�h�p KKS�rp�_�*0`��̬r���FX
��'JP͹@���X��* ��[�1���&�Y)&��!�!� @!"""�!�!�!�! �!�!�!"""��!�!�!�!j5p  5�5�5v5|5�5�5�3��3��3�39E9 ���	�H��
vf�	 AFFZX[R�Ѐ�r�
3��H  ��$ ���;�y�ȵ �����_����D�t [3�1�Fm�^���V�u�=�#�?�
9�; 
�u1[����X[�0N	P��R� �;�r�ѸM5�,�
�T5��62�6�ٵ,��%�lD�[SRy���D������c����A�XP �tu�F	@
�0�t���� ��G�q�( �`��&&�����" ��I��*.���qUFF-�+�R������n)�� h�QX<rI�3�.RS����Z�1X��[����*"s� [��� &��@D��XX'O�����H��$�I���鱲���w�[�$rt<�LWPq� & ��� �XRp��'�8� �%qt	c���S/�:���5@�pq�[� ����=
�P�c�P�P�/[qty�'��.⑒���4(L��@zђ���WR�����u�� �(Qt=s���#�H�4�I� t+B4B	Щ ��2����2�k8
eV����^1�Y�Ee;r	��N�	q�B����o1�EtXr�	���~  8
O���1PS��N�&�?@w�It)[�B1{�Ĝ{��v�.땸N2��&r����5I���2!I�8��1��$$���$�ڸ����'��4+���ؑ�AVW  �&1+��0H���~  t?�)��>�- t	��6�-�-�>�$eQ)u"`@"q��X�*��M��u\�P� ��{��
ԋ�p3���+���  �� ���u�� I��t���㣀����*���-��A���x��.�g�uB9�m{��p9�{t���(q� �h�>�]���,	��2���X��F�`-'ɇt�����`_^]�`��R�2䣹�B�r��)������GuX���V
0��-£��D� �e��9����`q� �[
�xQ,}�(�I.	\q��_qtNN�d �quⰉ��Ёq��t\�1�* M�+�QP�	��"��W��x͍V��������*�%�t$&�|t�@��p�o�&����f��q���랸�»��0��a�t�}]q t�= �ܡ���� �44�[ dt�� �.e g��t�&d�2���R<GG�X����t�Jv��PS�C@��p���� &؋�����}<5�; 2�����W��>.��<^��t�l� �y�dq���fq�ppa%$/���|u�=�*-P�R��R�	#I���"��c ��"���@��y	�U� ���:�tw�6�-���  �ǋ\�; ��*SQ< u2��fRWP3�`Hc��`$�uK�&` a��-3.q��-�,�Hq��-&�=SS�<��g-Q`q��u�B�[Y$�Z@wW2X18hX�t���1���� ���  tX�1�J��A>[���%���c��t�&%q���l�t� BG�6RP��#r3�R�|�p@t0m�9d��t,۟qvw#Qb.vS:j��ӥD�������&����H0��@����uS�A���t����S������	)t�Aɳ˃�0���� ze/3x,�% $�9+� ="�t�P�QPV)Yh��}��qQcY�q�cx��qge�G���x���8:Ɲu6�1��P�3�� ��`ϡ7�u �G��4σg�W$,<�:ĔdQ� �J��"���H��R��,�ωY���^��tQJnQY�BF�t@=�����8��AA��Q�A��t&5���"n��x`��@����?t+��ڣ��ҐZ�����Q��3Z  `��"�"�"�"## \###$#+#���(H=7�z� 3�@ZR��@��8����o�~ �������&.'7.�^�5�v�F�3� �#�(��� �y]�$=`7@uH��QAHOu>��!�͊_��q��b���3  �G��&��g1u��!
���;�����X#T�dt�ƀ��������\��h.I����T<�㻋�I��ŬbI�8���Br# �V���WQ��+ ����A����Yٰ�_^�o���qo��]��OQ�u����Yr��L��=����1�

������6{�(2u�_P nh4�4�4�4�4h�~���
�3  . � �   !  1   U  Q  R "33�KQQ*��6I�<<B�<HU<;�� ��n��4�#�������3c� !!����A���# �F vo�	����q������3��Y[[ !���qF��:��A#$'��X$ "Rq,,J��"
bl2<& �2+p552344
(  / :	,+8;@�+�6= )  ) (=A11+.00	,((>`*/6 9?)-�F'((
 /5?kwA";abcdc`eaat���9� fEp��>J-����W������e 23��_��N b��VW��2,��3��������������	 rˍ^� �(R-�u>ك� q �&�p���p����p���P0��-Ctd�-�p;���
���K@@��He��%�-���-s�G�� �����& P�e#����K�`���4��	�q l�78&�% n���.�� gI(� �?r��.��x�(-8��X��X�+r���Ƥ+X��2���t�;s� �� S�a\��>B	�����v	����Bʟ� O���81'X_^��]	�x��� �nVW��3��F�2��R-�^��^�ݡJ-HH�F��p�6���9���4��n�t<X�6q�>�  Q��-�� �u��t;�w�\ 0�4��;>� tN�] 0M�}����f��@�3�9��Hl�EXV6�e�K`��t� tḌ �t0�:�������)��r5R	 3��l���Z�g  ���p�X� ��� �s�1F1�E;6s��� �GP��؀��+ ����I��`��t�&��+ �k A�@t4HS��B�6`��)�%��HhH[�^�.;�v�����y ��%��5� �[y�A8��ðl�;e�<�u+� x�u#��u���m@u��\��3��� Z��R�@%a��p4�*���W��H��l&��6W� J-�l/��98���WN ��W�v�N 	Q��Q���|+��Y�6
W��W���&���^s_(m p ���YZ���&�oµ���ӲN8�Cưm���3l9d��.v;�
�����5�����v��ʍ7���e�����ے  ��% �����u�
d}�t}�.���M�t��&ĀtI6F�R�E����Q�˰�d��F�5��]�I�������� *��@r�L�=�s2�@ �+�� QRVQ�H�m��EZY�C0 �� }�����������Sfu�s}�6$�
����)
0$s%�&� ]$&��'�$�%'�'o$�%-'��'K$&��'�$�%0	'�'�$�%?'  �'�$�%�$�%�$�%�$�g%�$=%�&�$�%�p�$�%L&c&�#/%<&�#%0,&N'�#%4&�D"�#)$ c$$7$N%�&�$�1�&�$�& B9BK0T ��K
�u�|�:��q�t)� G�Y�j�>̠ 8NN�6lV�[w��i���\1���sF	������ ����X�� 7���I�Z�K�x�6�sL��&%	&����t�L��t�*����V����y�}z�0�: �>t��51ƽ��t�<�����/�������	 ~0�/���������=������tV2��9���=��.��%��d�`-s{U�辧�胻[u�� �[��P���̬x�3�/[��\3�6�{�6t�T�o
�_��yЩ (64w(Q�- -���'-3�
�P)V�=�Tp(���� ���4�聚� .<�)10���X��f��jU���w#M�c��	腀�r��4!�0�*��z!$� D � r,gHh�HS�����jyA}�;�X���S���1;�a$Fo+�c�ay4�&�����Pp�&��볮��� ȊG*��Xr�V��yb^_L�Cg2��=��J��=~�	2`���()�G 5���lJ`D��?��8�����U�\�t
���AH�� søD���y|�]��f�-8���u�PV؋GM8���B�?@<��DTO�2z�̼?u��0 ,t�^X�����	�#�Ǒ�>w� `J��tP�/�vX� �/ �n�F�*!�����Py�� �ْ��%��VPR��?��y�  B�@ +�ZX��
��t`�9F����#Qs
�u�f��� l���YA������-����  ��Y*��^�%&!#I�$������F�F@�f����H�1��>��D�G�x�"rDX���` a��6
�y$� 9.���{�F�7��%', �%�N���|���%VQ����t�*���6�J�scX�`��@A:^r$ |�΅	' �' ;6qr
�>s�
��#�&&�G�e�S.�����%Hu	����)�$�]c^[� �Hu�>" �:�����1B4tPx���C1+�+�1L���[11�٨0����q@�M�]�#�b��`ap��u�~ &q(�H�B<��IFFHH��� ��� ��Q��� 8@� ގT� ��	 �0t� �M�0�c�(�pn�4��� �f�#zl���l�p�+tϟ�%�xu�����3ǩ�f��pv+�GU�g���� H���u�o�q�9;�s�]�cf���P�N� �� �q�w���9u�D ����� �+4s� 2�s� �H��X"���8S��\�������
�t
^�|� �� �f`j�UCt����G�w~��f}p|#>~i- �* rw�F�6�b`P1�P+�6  3������;~�sV�\��*_��A4���Mg,u�^�9�*���G���ɋǈ�?+G��X}����OH� QP��^XY�nd8�� �L�=P��7� ��}�l�0͓[k��|
r��bj�r�;�s��@)rQ �c��[D �V�tI��W���VY��>������w�&D=TOtF �	�G��*�  ����� TGG�O ��l�~?OLR� z��a�^�쑨��`��<K���� ���IIQ��ي�``,�r&;^����Y��#��Br����Uc��T��� �'��(O��n�ȸ+�w�a�  x��� �O�H&�O�H !#V2����\����A
�t:�R	�x�;Sd��`�W�~�r_�^�  ��&uP��+WXt*``��	+��&�4  ��3ɻ
 A;�r3��� R��0�X���p�����P֒ �@;
� �&�GG�R��CZX0�u���+&G�� V���H��]��t �ˋ�I^� VjP��Z�? u wCH���<E���Dt<.���#t=0h*���
�H�\�ƪ<�� �u;�u9st �t�w�< t��< tN���^�W� ���m2��"��' @'���Q2������Y  S�[u��G�׊�_� �   � y � [ j � � I  �
���
+��06�� ���������f\��5���LE�a�b q "��
hʧ������(���r�t��<B��F�D ������ ��(8�~ /3P?8 <z(�\y<lz.1��)�  ��ncLT+4��e�` ������Á�3�-JTJ`4B
�V�c(��1(*CH�0?�� ����K�:4�!J_fH����nr,26/HY�L�JF�Xd3��4�DLlv�2j���`ND�w_�\fTep�v�|b�*��h ���S
��7e>�,�f�>wu���E
*�Xz�^�EO����q����}e "��� �l� * �% %qA�`HD6L,2�H�� )È (88�H#<+XH��HL&%H�($L= < > =>=<>-c �-PX	1 )H'o�>b_�w,Ȉ8	4gL�0D>K���D��s�^XX,̫A�
�J �Oo� #	��,L, ;r<!l 59Wjv|��E�o� ?����<VL�(9(*,$8,N,[,�,�,5�D0�48�0�-8�:<
�FU<bw��	DD$D(<D`DrHHJn HvH�H�HL'L/uP�D#TX)�$-X3P+ �/ = : (  .�=����� �����*4  KS[av
!-3�3�� &2�> T��,, ��,,,B,f,l,~`�0 0)0/050;�8<B<I�\<XDh}DH?<	�2H;�a�#H~H�H�H�:�82HL>P TTTT>=> \ �  <=<W�ی�2�"�D0* <>��Y4)8^ -@\PnH% ]�����?��kಂ^�
�/z� �V��.�9���	�1���%	HV �0���X	  ��$INCLUDE: '$ 0STATIC$DYNAM	 0�� �����2`�������:��\�>��%VWP���ǰ'���<�IX�����_^� �<3HH���@Z �/��X��S�e3ܙ
D� �YPH���X% Tk�2��,��l�$���?N��/ã*��53S�=���&����oCo���0���% j�L��	 ��0��`d������gES��-�!ӫ=`f-�����OFA8����l��	,�>��9 �"&�<�u��.#20��ݫ��t4#+Q�F"t���L����8bH��*��
8�Q����Yt<���k�7��@�)6\�&�3���P�3l!/��Xb�t	.���+��@�#	�����\ ��(I 8]����c�#�N�ff[�wҘ��31�5I�H�/3��&�$L�+�j� �l=���*R���<�}1�eB�'�l	+�	4�h� `$+���	��df�����*fvEY	K��2 �������)6���1���t�fRY�2��$�Cc��a *�=\ ����Ÿ =+��`��=�><T��� ��u����p���o_����f`�!e����������8�T!�N�!����r�,��j3P�i,7�0�^8��+�aR�H�7�n��'<`1kB�f�f�_+Q�Ᏺ� �9��5PQ�*���X�@%m
���	�_�*�8�!�Ә=���M���P�*�0��O��&�� m�<�:��0��@$�&��g�� ��2E`ŀ��t�;���v
t��
�!y�N�Â!H�u�`��iVm�!��ƕ���n��c�o(���1HdF��x�G41��U@uE���6_�V60m翎��pc;�  0� 38 D'-  XDAH[, !"$ ( 0 0
 	��@ VQ���.��4:�u���|. 0���s����Y^ÓfRJzCf ��	��7�T�Ñ��$� /�������a�����7�����`?:R����ff&	�	�	�ffL�����r�m�g�� T頙�	kY�锌d<	%r��� o ���t��8�蒹`��{P�o<�e\� 
d��B!�w����5������`3e����jH3�F��F�������)����A�̌��)
,��h��v	�X��q�8�"�"����/��A,�&-��dǁpf��[�����d&�B��Rn��$
H����c��ȰB���F�乎@�1�Za�(9��
1��K2�T��'�@H�)8 "A�\�x��3���"!���晙�!x�	n[����s,���rt�uj�
����
	03�"�.�3�	�M$��6�ff�30��f91�fv
�U�03���������	H����#�A �45�6n��	����F������GG��#G�+��Ù��{��v��
'� �&�ò��  �߲�ۀ̀��Բ��=�1��*7]3�N�5A����c�~X%�g��#p�a-u Z��p�G*�6���&P��TB�@tZHV�� ��^��XR�9�[�0+Ҁ�0r�9v���7�`���á9����V�/E6$�$��R3��'�w����1��F����G����l;[p�ð(��)j�� ��y��+�gd�덭�Go��|"X���sR��f��C� ������P�"��p��X��Q����n��iR2P252n�2�+Ɋa���>!�S�S6N!�6uX,���G��W�����<���� ��X���l��HW7�Z��,�? "���, �8� A5�HN�C���NC��������(1 u. �Fd�a���GR���
`�MSEM87
gfw. �GW< { k � Tm�pPq� ����<��.���� �NO3=
�k<̀>t 
��"s�����O � # �2��3���fJ �$�~-@n����"�l��$W,:�P��� �3<�=ùO45  � �!@��E���� 9��
�E
�(
H	�0���d�/Dx%�/����&���H%xH�@G��r�3�A(�ʋܛ6�7/6	���FV�I�������B��0�+�������! B����PUN���v ��S�>���F2���u
�[���� �����u�@�3����E ''���  ��������"�?P��F-�=�� t��%8= Xx`u4y��n 	��[�]���X,�S��6�G[ X��VSQRW�^ N�ӊ̀�8� ��˄�tR�V0�����u �� n�@u��4`����tt	�'�    ��?�6 ;6!�����?É���<��K���J�K�Z=:5���Q�� �+���DD�f��@�@,L:�Z�ZQ��uP������%>J��}�y.��@�-21<t#O�VR�U�V=U��8��F  F��ʀ���P��y��{���a f����$u$���{�_��n��À��Ff  �_ZY[^�g�$��
0��� Q�Nr�9�8��t2�00uT��V����V0;Q< ������ �T Y�N�M=�HM$��^��9� �1m�h�� f0$�@Bd8ɛ���،>d
Y$��B� �~�<���t �!�F�u��n��~���>@"3�3�p3C��  �%���=� �Xs���x��@uOWVQS ���ـ���؀���G��#� ����v
��V�~R�s�F~V M��^[Y^_�00�S��Yu8��`u1����+��0u$������  ����u���u��������� D ��   2 u��L�!�[�s���u�.�f����Xϣ %<�q0&��.f
�
��Õ���$3�?]1�"7�% 8 5�@>2������u�G��LQ
�& � U�2]��gU�E)IgE�
���N��]��� E(#�$�i3�	� ��N�.���C?"G
� ! d�tّ�z����P� )�3P`�� -  P�2\��
�
�
C�
<x�
��
�
����
�
��
�
��_
��
�
�=��
˴ ��������{�7  AK���W��  �Zc:��n`>�(G  Nu���������!"7!c!
f�"|�D�U���~H	$��/C3�{A�)x/��J�^h'% hk_ Yc:� 0@B�,� [�� P��@ �y�@���?���}����R8C6�`��j���0��� �Se�B׳�#,`�k��
�8�d����3��9@� A5�h!����� �Kx����\)D�;��D������ �\�y���r��P��{Z�>\i�<�7M�,����2Ӏ�f�ˑX^8y����2 � y�	cf���p�9���F�����2 2[��ɤP��r����Kx������+�RJ�+ l eBPU��<@��K�$��C�@p�8V
Ob� @c�m�QP��;$m[ �P�u 2Z���t����T=��H�_��J���<&ow{8���
]��{����~�	��-�~w��� Wq�:�O1�5x�^���K�z��Ӳ� ��(	/�>�ĊX�@ vp>[��R`@�3���&���l ��_�8UV�� ��vNN����^ p]�q
|
v
�
�PܪRQS�� ��Ӌ��~GG�`�M������2��~=
 0�F�
�ێ����P��F� @P>�؎�BA0��4����D�	�D�)��H3�v� QB���@���G�,]��?���K�ƋV��Kԉh��9�%  ��Qp]r���  S�� [�������>� �G��@q�BߎǣF^C9��z AA��l�H r,�<�63".�<��F(��O�&�Qa��a�)�2�+�9h�!�� �Հ������2�+�;>�8����]H�[YZ^_�g�8�Њ&���D�?
� ���e`	������T�`�A�
 ����"�*��"U
������s��$��
u�@��t�����TX;�uk��F��=  t<�(A�����MGij`(�8x�"�R��� �\�t3��R0 6@ú���� �3`0һ������	��,p��ZE��
D�v 	�2u
2T
�8M�D	'����@��Q �U
�U�2 �=��2����� ��[��sR�
�(���.�ǃFT��;�t����2�x�놴߹� �w����`��+�|���� �=C ~/UR�u���4y�݋��] 1}J�x�I��00�� ��� �/fQ*��譋���ح3���7`0p��|5t�ʴ���zu���w�tSr)��|3�W���Ċ� �֊�͊�ߊ�2`�+wt(�����`����Fu�����?5\��  I���������΋�����?�X  x"L\|s�/��,�,s f @���}+"� ""����������������� '��X��P  �U��2�R�@P"�3��ۋ�� ����t����U��U	 l�ڃ� �D�&*XPU�P3�2�����2��Ik>II��I�I
�eЬ�ʃ�CV{ZVգK0VՁ��?\#O�\�RM�=^ӫz����Q�DU}����� ��Y]���a3 	�^�a ���2�URVW����H����_^���}������ �3��r����  ��EU�> �J �W;�@
�<8 ����c��r"�>;Tu ;�u;\u;s�����
����Y[v�<�6� f;�sb�u;� �wA��RS�3���Fĺ���P��aD���衚3�� ��  [+��[�]蕒��scO?7�.es��O+�{ o�@��ɰp��u^��׏����?Ո��AUX]������ %X��  ��Ǌ��݊�Ί򗕊�C�2��!�ufNMDs� 't��S��
��tD� мk�r���wr'� �t"�XP��r�܌���1��*Fx՚��� � &p]s��
�
��~������4�d�–d,��t'R�dd4dX��ݪ��i2��G#׫MAM��NM�Mk�M�� � 0��M�]�EX]� ��e
�� @}�~`�u�E����o�`�����rwF"��B�R
��=�Āu���<6t��p'�&����Ѐ���$�ȆĞ�������ʀ2�  �!< t3�d
,��D ��t�T�|�x��D�D���9�����q�-؀���=��ɢ��I@H�瀋��
�y��\�au��E ~u�\�D��?����� ��� �ؘD[a sD
�L
�u�
 �=� }�=��~��.�&�.�<�T
���T
t7���<��cr,2�� 0�rw��t�Ѓ    2�y	������t����ë�,�
�x�돨����M(ՃM1.�
� �
�.��8��ॎ�lF�  � "����M0�H����=�7�����
ƋT�87���-�s	������L $oފ�2��%� CHP�%
���p�҇��so/�Ȼ�3"=� �ˀ�\�L�T�l �ʊ��t
2�&,�4x�m=�t=2�-��h"�� @���u����&���3�2�,��L�c	~�y���,{��4r�'	ߏ@��)�=96AD�L���ګ �� ��«�|
�瀸��`��B� �\p�����L�
��4�V�	�Vl}߀/�~܊o�$����Rl�K�:70t9tu�4�������T�� ^y&EY|�S����s��:
r��N4�@.�����
� 5�
�Ã2���-���P$���q�
���
�
C'��	t��R��0��^K�̓���!�IT��D�l���_�ݐ���Ԑ�T�gl��9Ӹ R�u�2ɀˈL�π倀V߈l
�Y(U$M(3��]c�8eD�O����V0�Du8`u.�L��*�s��|�`N��*� �!
�y��t3�x	_�.�F�+�(ds��8��t=������	L��������{����� �-,�V� �m5K��A�2h�3�|��u!�`�]���`� 3�x0���������M!�Ú���#�t?��?���sr���~�uu�����1R- ��r���@ ��_��@S��O*E�5�?A;�º �E^3��x�ҕ��H�3���� ����u���\��q� �"���t��HsZvj�} jP)=����K�-"B2Ʃ��3��������r�������B���3�L�W��W���?��I|at+o@}[6 �~��t�׻���$0�9P�Bs�������u&,\^Cu)u1
�_�"���s`  ����ð2�9PX��)��D
�u�����]�Ͼ:�����ڎ�\؂�k&���;i��m�2�=�A�%-�?�q��|=du�O@0l,u�[���0���r&3�l�'#��h|�h�`
櫩!|�����l��]}$�$ȬHu��]�!a!X���~K�|
D��u��K�g4-4��d
��	5#m�ʅm��&�R�� !��E$ 8*ȋE��M

�e���wp=�%=~?�y	�8>S��$\� ���3��.�t��e
3ۊ\��
]H �2�xF
�y{���;u|�Ybkhr	f�we�@�7_9Fd]A�+=8m�$�x�.��@n�x����Wet��ܵ��U�6�!�A\.Tq	>���� ��.ע��b�d2�h `t������a����� �B�,�
��㩋�>.�I��`�sZ�����%1�!��������F�[t���.�� �����FF7I�<�iU��v��v9���YI�t�v-f� 8(�B�i����Ua��3���~��� j�E+D�� ܨE}  ��B�;Dr%w;  \rw;Lrw;rÌ� �>3 ��!e��� c�Z�s��Qt\�}
(P�Ń���.�& ���N#���.��^5�b!ѝ�@�D� �~��3��a�W�,(�<@'�'�!��x݅����ód` ����râ6� �LB��Ep�,��s ��r�.�s���	���&r��8N��Ӂ-�DD
��u�m�V�J �EG�	�HB���T>.	@��*��  E���r��9R�u���  ��W�s�����3���\d��E���o
��.ȃ���{�]�v;Mm ��_`p���쾃����3���W��B��_�:�@��V�Ɏً0 9&�U�:�uEV� W	�� ��ʀ���:�u(
�w�s�����?/�;�u��Ƨu0`6�� Zÿ|���WVS�p� �� �^.��_R��QV���V�V��CY���^5���|@.[W���f�-E�Y1�Q3>���;;��;�_h� V*&��r��^�4�xû��]��'�D
�݆D"T%��$%xj� 7�88��s6�c��D���� C�,`����5�W/��@�@�P7�	��+�X��Q	�P(Z5�����$�H��W��'�� ����E:������V�X7E�1Ñ�d
;
]���D �\u��wH$#CS�����czm[_S�i [� h�t9��y0����۹PI��s�W��~J�IH!�O!c�d�u:A�N�
�rަW �J��V�h�R���^����T	���Ar^��î -�5�!�"#�`$#�Q#%�PR
.�Z X�.�> #Q� �� Y.��t����.�c�.$ ��� 8��v�z�.��0�o 	�^�s�d
 P�'O�]� +� ��N��eT!dxL���\���!Vp����v�P� �"+�3ct��! 9t�@u�3۹��w� w�
 �@��0�#���  ����&f++Ƌ�ݸ�3ɊE+���Πg+����+��,�3Ҋ0�"�⤠%+���ȸ��$+c��&(+^�8��t���UD��##��3[��u'���:+ u?���Q���	t��P2�H��2� <�F8&_#���������Q����5��>33�� 4/�m�^S��  ���OD�WFu���@�3�/[�َ��WaJ���A�VW�B�nԋ6!gı#_^�O�����V# !�P�=�؉`�&+�p X������ �Vo�

L
ͼ

B

9
8?
�`
. ��*� 7<s�(+�Hbku��-� � 0��RP��	�.Zj hË����%+��5�D�bZN2+`�0+�>/At�+غ:�hR*W+�W�,����u�`3�����a:&8�ؖt@C�!�*��39�4+2���r��_O�Ί|* o�PPQQ����N�>�o�$S�T� �!��A�.`�"�&;�	
""���B�͊DM+��ډ>�@����   ���>
t)�]+;Ā;*r�^����G�`��a�+�]�R u��WV�v�~ 0�l+�E�ȈF�� �*�F��Ɗ�P�	��E
��	�&)��D�m���30�	3����a>(��a�azc�N8s>���?�V�%4�Ft����~��L���- � �/F�J�vG����kZG�D.o]JN����!�r/!!N!<� ���s�R�z`)2�*�+�-?�!a~e�9��
s�yU�N�$+��i� �1?x�MHdH9�  k�$�/#���4I��&Z�8":	^_2� � ��88�>D�fn`@@�f+w;~�wUn��g+G����&~�'��T��#�^�W�Fr�6K舼U�JPW�i��P:f
���^
 *�������
F�LN���V� ���׺^�+��% �/�
^ӉR62gx2���K	7���s2��d6��F�0a��>�+�����-� ����>�- r/�qw'��j� r
wi�u�
��
+������������*���������J�x�ZB��l���F[����v� ֋T9Ww��pr9G
siv�&�rnrKO��6��� ��� `���P�� ��������$���"t� ��6.,�X�bH=G��a�[�i�-R�&a��@aDa� �"'��e&��כJi�'�=6�6X�f � �;�>���أ�0B�k��;$� � rwS�����A%�}� GuvBIe��Jc���ވLs���7���	(��u�����v 7a
 �
��剂?V�
D*�<4�1 u' ��-t)��|u�C � �u��~� u
`�6���yu�*9��a�v�s*��A��u?�:�X=S�;�N8��<n-�F
�u�%9wu ��1�=���W�y-a�~
E�Dv��=�=~���w�;��v
��rz��qh�!����|�!��>LF�n��&+��u<��~8�u	���	�tT	�����13)�����~���.z9'[�m���`���V�6(0*/� H��^�?8�G��F���G�σ5��Σ��s��?FO:)$��V
�V�C	GWԠ$W& �8D�v�Dw�vw�D4`%:��	�t�
�uԛ^:L�o�8FT�,!�V��q����>H�� �  �z���|=�*�<�6<��� �(P�w�q�%���y_��C���E�#u�)B�<�&E�f�)			���w
w�L~� 	T�@��b���-�Y�ġ6+�8+9u9��t!գ�����
� ���� �|��u>�t-)�h+  !��+�;�wr;�spB�DF��$�B�R-뱍MEEC�]E��EE���EE���!�-�f�^�1�h(�����F� �� ��˃>�68J*Erx��w�|ot�>& �V�F�F$��� b����� s3^��HM��=&�� 8P�4"4V� W2(FtK�N�G
*NtC2���� ��^�� �2�����J+���91�< \QRW�� _ZY� &>h+�Nu��/j1_^��`
N�xN�L�O�z vP��OK
U�::
+:�v�r�P:@:��: ����Jw�q�US���6ohQWd`8+�4!�[����s:�u���
��
�u3�Y�1h�#���2�+������.`M�WQ��X�SX8X]��l��+`�2G�����u<!�g�T�dt	��[ì�݊�����>��� �����t��u	�p��		t�=�����,	p	*�ê�G����i�Xڣ-+�GZ�á^�/ r0�����P3���  3���p�g+��RSP�x��׻�P��$! !��.�?,0.O�(`!.4:�d����؅D9D�u$SU��^[`�T ^�L�L�Q����+��^vgcK
�?tx0H�t%�d���?�L��Rd7^p�VW�:+� e	��� ���%��O�p��� �![8�G��2���h�G��,$`�j+�*@�7�>�Jr�D�F:w
�q*X��Fr�A��We8�?���I�{�!�������o+��� u(�2o�"bNWPG��vV��YX�@��_�\pE��E��;�}SHf��~�H�������e� �02��������p�[ ����tP���&��
˫�P\!�)�����>�N��8!*E�H�H�iE��QR+PR�6������ZXP3���Hu��xg�Ot!��Q�"^K.� IL�p�G���O�5#�}���� `��9Fu�.]F���d-������O�sN���N(.��4j��G�  P��������&����6\sa�q|���@P�X#�� ^cQ6��!�W\NP�Q�\hMP<���U2�+� t�w�����Dv�tL���o�G�� (9?v�S tҸ�К���Ǻgu�����Y����t ���PQ\��Σ<]�s�J��Ȫ� ʈ]
� s3���V��&6w�ڇ�����ܱ.2U�|L�u� �~��v
e���>F!~�v���3��7�ɓ��c$�]��t$. rDt]FōB6,6��Гft� &�4��+Ҝ����(�Jܹ�.T �!�'���� �#�$�X�H��£���ŗ:a0V�\�|�:����,����-' �
���O�-�z�SII;�v*M�(xT+,(Es�c7��� �E���eR$$}��-�d���+	@@����n�$�>B|�2 ���P��]��-��-E�-~�\� `� � �lci�]�@���8�e�⠌������,��-�>#!�Du
S�Ȱ��� ���*2z�� �M>��JrJ�\P ������V��6N����rG�	:�#����pr�tQ���H�M��AD�k�2k� ��ma��u�W��n�Z��:TI��E����HPV�|��ӌ#�T}�N��J�@I/�m%r�tf����
/%�K�-A�����6�-�-�?}�
^^��@ q��+����7+�� ����A�D��
��JyUEh�� �ODqBYY�Z�]33�/�$`���T���@[:�����t��9�t�N8L�z�uT%��Z������_%�w�> ��t9V�,����gP�{���GJwbeJ6^�������u��!f�����V���4y����
&1���d���3/��?d��n���ڔ�!g$\����w9s����\������|�-v�����&a]>rϯㄜ�[��X�X�X#aT�s$`1;7���w�N�D��;�rX�X�%?N(V����U�b�D)F�<[u~�q�q	`ƀ= t	Gw�		u����H�P��
)�� �L)3�F$k +A��@%-1@�Z��/tu�
S�WP�� ˈ�M�v#GW�p2S�F+H*�)Wu������G�w%�������	�R^����@����v9M+�ր�Q�'Kvr"s��XXg%��q�������C2o	�@.L:5@��0R��R��jx�Rͺ��d���eG�4�t�O9Gw=��u	�Ʃ�I�  ��H��������p�v�@�0��N�N��D�A�����^I_�V�����D0�*�E���!@�W�a�]��m�؊8:�����P+���ۆ̽G�q� �2v!�ƣ�qW��Ƌ7f~�T��s\���#At�&�r}���?�*��6��wш[����A�%.{�`�lڀ�p�F�ψh�/ gG?kt!���HQk����?Ȑ_��I���;X���Ȁ��/̃D-B8Fv%+!U������q�sX8>rXs����d�c��8���+����(V�����x� s�P
��v
F�ɴ<tFYA��:Gs����J����A�e	��8;V녾����	*Q*�h fK�)���om�m�G�S=$v	.�tIpc"�D������'�;�tԡ	��}�5j��1 7�öDr��6tAac�}�pN��f�>���Ki1�@ M��������t�u�.q�6�y� �ۀ������L�F0�u(F�1!�>:��+����1������ ���|6�r_�*��4W yW�"�$����Ua
�0Q�
b�~�c�Y}�"�8��D�K9��^�G/@��x�	�ǀ�	2�e��&H�-��i���2
bMHI�@c���-���Az�A����V��UB�����*]tf�!I���D=j�=����=%*/='a*.=p��p� �l!Z�=&)R� (J��4��nN��Wp~NQ�tVrM���;����K5���=� Ԭ��a�N�p�z)�6� o�_����9�W赍���(�Dō��<�'�tϩ(�t#���Jk�T��p�q����i����Ι��N���v0�� �����M�mG����h��v���P���f�I��� :sw�ovOud! ���P�Mg�=�@����*��PCd-
�@���^��x*�.����9(�߃��B#����%�Eb8�� Varzw�n� N�c���= ��vV�y$�a|z$T�$$���$6+���vk
A�je����K�X�c�L$�N[��v?��뇣:��i�����p�^��7S�&6�!�K�e����� �F��x�d�,ML������9j<x3�Q�fm55�1�SS11�J?d��533
�@��%@m�-e����]Gu��k��<ɀ��>���+x�Gt'q���uNY$�� �j�Fg �@WV�NF t��F��W�ݲ�p��-m�������)��Q�X��yD�މ^芏�!�`�ȉN�`A�A����1�<�,)�4�lf&;HFF�v�����9|K��2���7���F�;�wȻ�?+ � ��D�=��P衾�t��� �P�&��Ƶ#�"ˁN�����	�"�~��g�^-��^F���lB�tuWd Q�t��\G���p�_�>p�.뜥8�&&ǊN�?1>v)M~��9�Pe�H�'�+���A�{���SZ@FU\�O������2�B�݆��Ƈ��q4��Y���<!��� ;�f��!�X�?�EA\�E��~\��E���Wr����WbL�s��S(���n����'	z����;zM���`�6�p��3�vL=��t=�tR=�X��3铏>�d/F�0�
����Ӥ{&a�V�I,&��i��w���Մɕ
��u<�F
r>Q4쓀�'N��
!K~�����98�`��� ~q�ȹ
�;�g���xP�F��-��ӧ�	sm�~]�;C�!��-�N�G�޹~�-Q�-����-8s7��s �(���R�P@/� �~ R ��ڤ( u�XK���P&��eo�w�{��U�P�'������X�ɨ��@Cq]�������<�sW�j�]�-��kO`qF��^_m'��4�W��j��f>��;�tlW�<���9uGxtV�@k����^��vT�����LE�&Y��  ޡrr�tr �
�V�H	�g	�p����\�vr�4lvG���> u�	��[H�pO�O�Dn h�fCm���2�Y�q��X蚙�� �ƀ Ł����D,�m��4p�p �|b}g ��8Eu�
iP#�	6V�v�Dl��[uK�H-��*(|h� ��r�)�d�F�~��~~Wm�B|��~�~p���tw��A�є������}�ޣ,,>����c���$P 
���\.Lq����(A� �e9 t �2t	�2ԁ�97tz���o�~�%s	���><)uH���B���'��u5(.�\��P�u$�F� t
q��V��� Q���@� �� ���ǐ�	Ʊ��� ���\2��D�H˸� J^�;�H u+��9u
ju�u��O�=���0O��vB�B*�=	�ع"\p���.p �֡  u�W��w���rr����V��' �% 8= uq�3?t	�$?<	3=G� ��W�	h�Y!t�C��������P;��F��g���p+ۋ��jp�})��OhQ�~tw�<h#��R(�>t��r� �|9��h�1;���09j����D&�W&�����x�͇���E��
������ϠQx�[�Aƃ����Wsees�tHju0��d{�`���l��5^�V ����D�ˈ��VU�&D*zW�Wr���W(�lG��}Z)m�
 ���9 \i��E�Nѱ@H�\��u%*[�T]n�(���'u�� ���͆ ��<ar)<zw%�n� �2w�"%,��yx�0rsDZ<�j� �61��v��W�m�)`� �w',Ի�� )�� �� ��8ukp#��t� �� t�D?�~|�~�L�~�r�9KW��u�y+xX��2`2��22\FIB�{ g9VŖU�U���t"�bIؓ  ܀t�V���xh���9xu��[ә�k�GS�.��"9�V�8�?�՚�m�c�>3�`t�N�7��d�]��	��4(��_�5'Z�PW�r���YXQ�|�ޅ�VW��,f�����TM�^���4��%�Ȋ�+�AA��T�s*�+�@���-^�v�
$8Fr2L2s}��5T��O�(1sd}�a
��N+��A/^���~���:s/G:E����1Gs��EG!�GV��0�� ����B��x+��_�0/�g0c� 0pv�U�`��W�JWK
���T�
M��v�/u�s�GO���v�?�����z�Gs�å/09y3-�r!6�%�@}U|+�e�0�X+ �GF�dK�V���1�j�*oF�k?ޱh�x��@ U( ���=\1�7�.11�1���1�1  �N�1�I�1t��h.=��= aD�=d�� *�DB� !�<��a��N��mN�0w6�%��?
BR,�O<V��`t��5f<�vנ�Ln�~��T���:<��<9�'�<i*V9�*��]��=��  V��'  ���z+
�
x+�Y�.�8\~�R���s)'bv*�F�	\v�����<�hXe�Ƌ�{&:^��* ��v+��96�u�PG��F
�-���^#����ߔ�>6�-�Td���>��u����ns�w[2�Eh�| o5>t�sWZ��# @�� }C_9,}��x,;Gt��v�V�D�.��΋�+�>ɋ������&A�V"+~d�V��'\�=/#�=v0���>rw�(�A+������3��l��&a��rHV�A֣�\������To�t6�@i�V��&A#R��yizj��%M����ݓ�k"��� �V�^����1D�0��4G���dG�$1�S��^��S7
�/T.%S���B?��t �C���D�����z�(���K�t�s � t���M�w� '��T�I*c �$���밚X�%�k�Lw4�~�-�!��R�-:��-Q� �.1�-��!�Ív�$�!�+�6�X@ݞ�xTƚ��-��]-g(�N½� �L�f���X��6|+� ���5��c @��W�D�T�L�e��M���L?��Ɨdg2 �T�F� .�0bF�H���~���E��q�n��5��p��tw���E�@<�@$��G7�t9n��l���Jh%?�N�� "=0 r�u� {����ʀ�ˁ�;�1�A�����F�l.b�	���U��0�	��&X�s���9��-�|$7n�|�����-ˏe-�#0,�
������ ��@E $�����|s(V7�-P��L*�����-'"ǘ�Dm,�����S�2�yV��KB.��C��B�F�t�b���>�i�̎���p�(�Et���	����!�������l�;��K�~�Vn��؝U΄�[
�f$��ή���Қ&���Nؘ�u4(���n��GB�@rĀg����		��lxtҪ��4��\�2E���%O?�R����G��t�ڃ�&X���Ίƹ�=rΣ�=�	@���Ҁ 3O@�G�G	�_ ����a�]�����}�^s�ւ։�0���}h?��t^_�*� �N���8.xprt�����"�<"�	8��*�N�"T�����<U�0�_`;9J&�<�?��-;���� '�.���;��xCԀ�?�	�� �r�p��Gs�
�Ita�����\!w=�*q�0�A���F����� �!�n@z�O��]����=ʀ� ��t�OS:v:E�9�!�d��/L�/�G0	 2[�4Ӫu5�`t7�?��_�A�Wx��W�rR� V~`VN�S�����f�`��U��XF��~�1�!b��`�m�wRx{r��!�O���� �3��F�U�j	���?0��0�6$�D6�C��8��9g:[:�9�: �:6;�;};�F��N�-/@�v^�u�r �u�*`/���V�`NO��q��D
�L�/�$1,���f���\^�ē>Xg2�A$sX�'�f�*�a�:GV(n��MM�0^��d�K`�K~���A�A��:�E+U��>��M����6�-�]�~� t���E�N`�u#�GH	N�D�&ey&C|������ �G���GG_1s�������~s��N��>� 1U�"�"|I	���L��{� �8p\�=A�*�-=
-L\��=T��UKV�_�������YU�v5�s��["�"��dp�D���&����(�� �WV�>�-i� @)�)6/q������B�b�k��C��u���^�gq�	�-��"��u�F��E�B� ��6buœ�ٸ�T���O�4�x�V�܀낪�-/�L�d:�P��uK�.%ny��쀆9��F�$�R�[-{eg�H9��*���+� !���!>��YZf.�ɬ �\�1G��V�� 9���x�q�aNZ=�������^+F�BBu&J����"�D��a�^f/4p�oyw12��ܚ���v��4����-/D�E%�=����*��哞$7M�����&Z�=� W�K��ݔ?��9��)s�z�	��������4�Q��4�&z�K�Xr�����u�����֠ h'\� �a8��PG
� oN���b�_�� ��!�!y�ݻ�Gu\�GF�(#�wS\'?�"&�S�w���I<���D;��M� �M��:�nt���PO?Ǌޙ�T]$�/����+�tF�,镺/�2��4R
:���X=����YwC�"D=���=���=+����*��R�a(BQ���@ �'��n׫<�	��� f��g	Mst�v��o̢	<���;t;�Ov_�>i%*Eu��m �Ch�!��K����넇DAv{���(�(SFB-���� �Ƒd�{G�J1�8��Qm��!��������N3�'NO	�Z�T���>*�����	�ႀ�$
�{I2,�	$� �,t�7�v3A���������@��t�Uؿ'�37����)E�.1t�R��9|� ���/���!����d�5FM"����h
v-�^��V ٭r�cs&pW���� ���� �����f&g9F��1���Nжb�^Ap��v��W�)F�~x<�\t/t:��u�*�~?�+���$�ΛD]�Z�Z��� A\.%�� (n� �t���~�5_U�ډ�S�$w�Lf�D
"j�DȆV|�D�t����5Q
�O#�"]�
1_�G Ge=��P^%[��5G�2��S�B�բ�^���H�&�n!��Z� *��BV������4��u�  vA��u��Xh/�_"Tb�F�8�����4�Q׸�$�UA	M��?u�ʴ�p�	hNP�G�t�x�'*R��i��,�����J��WOGZt�PCE!xGH�P���|'A`A�O70 ��RJD�N��
����C�LI�W��ቇQ�2�4k��E�"7��{�7�M��Pd�L�� |�=��`���p� ������7f�FLp�� 8GG�x�B�LRKs�^�7>�F*�3�f^�7s�F�Y~�Dm�S��^���j k4p
���_�@M>RY��H%�y	������=y�I�J��i �9m7�f!S���3����E�< t)�4.�S+��]��P8�CW����7@�K>|�������"9�`�؉�5)�rAd��G�]*e�bq�q!vӛ�JSD(B@H�Z"P���U�T��Z�PY77D���A6;�s���8	�@����S�D�Du���kg���mZY����
�F�!�P��F�f��1s$��.�6�|W@����v��PRW��cNCt'����sJu"4���o�(��6�Q8
��_TĴ����|`����,�k�@P��L"��8^S�d��	:�|���P�\���ԣ|�
�N�5R�.tEI�$�H�CuUQ�UʊRU���=eH�Eo�ڝD�~,�%'*N�DOU��z�g��G��fQ�:���V� �5�������#!�6H��'m!���"'�?������Ǣ�b��;��|�}��D�rAt t�V�R�z5�G������z!(TV!&2��\��&_�&�d��	�/"����sbx��,	c��Z���W�_H���ٸE��M�6�k�Y� �S�m�|.�dD"���UF�`nC� ��r�Y�k�.���!�="9),=P8�I�i���0�.��\�\f��IB�p��vdḆJ�P�n)\j���E��u��e�w	�D� �sF
9J��;�/��V�
�3�y*�#`	��!�%'^fA�]�N�.�4W�uy]A>�d�G��D/K�v�H΋L6A�����f��E�7D Ta���`z�~���'9~�u"�Ҩ
8����� R���XM'<z�O�	�7 �8F�sV�^
���)r��:�7q�+� ��rER�
���9|"}<Ji&��"�i�;�p�L40�"8r'�v��	{ca�H���v��w��$p^�w�V�� D4��J�}��"�%+,vA��	�j

D_��T��/��\s �Ʌ���ã��
B
5+N�a8�e�
���5�8k�-����C�{	����-���N�Far��������+D��^({��|'|�+�!E������w� |�@���+��v��#0�{��/HG���.�k
���V2Q���\�"mmTA�I��<90)�/�h���?�f���8�џ�
@�oD6�D1����0�؊D���G���G�Dq�!�9%�O��?S���3]J��=��t��{3�!8�_=�� l�l�y� ��I��G�=#tWw��e= Y!�D="u{&Bf2����A�i	�pD�P�.� �!� �X���AQ�2���" ��Ve�� =$`�=%!�r�=&��='�(�(��<�̼�ip���|
 r4������(=&�(�@g��d��?��{�ϭ��&�C���7�w"&B�n@�=A4B;��&��=D
>E�hHF3"DG��=H�I����	����&VnK�
�  ���^���c����{�� V�m� P
$m��tqN��t2:���HC�RN�	�G�� +�4�y�K��P�� vo+���}�Z� -|(.�)5RU=�V4ȋ
&�lx�$�s���l+h8�M���]��g85����%&�W(f���~�&&T�$���β���ɋM^
7��$��G�!���(�?78�;D6u�A�Z���7�@(7�ZՄh̺�9#t��&�a�(��	��-�W�F�L�`��66"u5�|�/]� �;}M:f��2��P�]=�=�"����K N����a �l�O��= �b� 2[�趺Eb�R2�H"�
�{\8�p��������|��8��
tY��`"�:��P�
����	�H���}֧<8$��09r�$+@��B}%�?BxBj"%s�:#�����v]��-CU��*7�F�T�P��	�P�h������6#�������p��VWF0H�����d��e�vPe�H�i���d-`ռh}Y&_��f�{zf2� 룽t;M�������vE�t՗!F�p�%����\���H����2�0@#*��"^��2r�%�w2T��H�C�C���+t
��/P���t���� [S�4�|"��7uW'=9H|w&�.Ad8);�w) �L +ȉN�;Ϝ�s�!��pz/�>� �A���*��@���qB =��Dp�d�vx�H��f�R�JBG%�z8��T,-H�y
��9wY�)D&V���+f�1;�;�V�S���L6���
��qz��� @J���n�E	Qa*d�b�]2S��0����� c_SAI�uz��!����s�[7�K,�eC�bD�U( �B@;D sL5͌L�;u4�Q����h,�^{�?f9D%"A���ALAd��A%�:�A��^,���2et������*�f����s�]�V5��2������Hi0H,��&�H�"��$M�P�¤V ���JT�s�6  +�|� v�n��)"�G9|A+���q&��Bdnqq��
5a|Zz��n �|vc�����A�'�{"�����^��&=���|c�!PdLJ��%VW��s��=b]޼���	b�68��C�&��*<0r���!<�
<��n� �f�����_A�8F?b蒓����j�ڸI�Z�����8 u�m��D8gW&_.��0���}�t�t$3;% $=利D 8�.&�^�*Vx J����D�\[q/ �IuH�|�d ���H��7:ǒ H������+���&����0��/�~�EHڕ�~�xY|Ø��5;�-L��t'�� �	t
�"/�!@��V�d
�*� �.�,�D&%� ��u/�` �U$� NF��,��(T6�*S,0
" $R�u�d(5�W/M�8r�,�r%0��+����"�jt��_�دtǃ&���$-(]0�;^~r&�*3 }b4��D�^��u�:��N� @��V���AN�<��d-�;��Mѵ������\ �t �n�&����Gy�r�&J�O�^�g?>Ihau��,$P�TRwK����S-I�$�!w|\$NrV2�4Y���֢2�4v�7ě�+��l}fF��r������mI Dե��T4��(�3���&S,�)f�#��VLh��t)�_�R�v��q�,d��L �(d����n;���C��rb�3�H��		��VGc�&�U�5{v$�c�,D�;�9D"rMR{�@�C�S*5��[-[^��*S U�B&����� �R�S��A�x}s+�����}^�`}vQR���2�h�+ς'9�cV���9"u%I��O��a�=J\O���Ф��pw@���Ҥ�N�e�g�
sF���z*�R1�K��V������\"�̲��3��;"����2< �]�v�记�*G�;�$~<.y�ز��)�����.��\/���9i�ѝ��@����W�R^	�G��K�������)��5���U�A��ja�.�Z���C��Q���5�rҏV
�a�~ŉD�[�	�EG��"��G�G
���G��K���D	���_?T^k�o�	 � V��!B��QB� �VW�� t�~��u	�� V��F�k�*���F�e �K�� �G�� 3��f�*��� 	�		������� �� 6�$�W
�� �� ���=� �ỵ���� ��w�� �� �w��6~ ;s�	q�		�0	�6� �A(}x��r��H��{�� v9c<�� �2 u�&���(
�[;�P�������Ρ:��0�  ����=E���D��R��e�;U��W7pI`K@$���	V t[#<w�z�3�sYDq��s3rsNs�N
"��4����Y��fZ�^��go"�� 5;��r�+���.2�7'IPHCLd��&��-'"�Gq�>�~��Ař5�*�\w��="��� �-w.�K;�v�#���S�FN���&BVWP�&�� �GMt5�F�� �^�N�V�PSQR���9u�[�&Nꨑ)Q[�3��Ĕ��gf������[3���=�C��i� �z|�)�6�D��0+"6s��%AqlF_��"n���	�ѻu9�{���N�| �t;�tJ���B7�@0U?��T���Ou
�� �� �� �	���YY.���t萀[	�p�	1�~>��^�x~�rr*߀9��Q���I�C@8�L<n�3#�ة�	��5`�% ��y�
��-w4�i�S��E�\Xv�/ a$��D��e!�&�9.�f�#g�A%�l��;�w���H�Ǟ�� ����� �at�{�dD�u� ��I�KZl���Gtޤ��&4M�|�!�H�#���
���r���$�4��S�6e���;�v`�t\	�	 ��Y��� 9����2��Ay�IN�w�z��5��  ��N����y3���ˏJ�v��յ���9��ˋء��؀S�_[��I��xN��Hy��/����'wueq�
� �a��堙`$g�m��۝;��}$�e��$׹���� 3�3��Ž��g���^�6� 6Ń� |;�}� �,|	;�}@��$?�QZuqf��� ��t��@tV�v�� L�t ���tp�� �r�����l�va�o�N�}(��0�SQ�9�M�w��y+�+��D#s7�#�z�^�*�N��h�fu(AniI9a'Ҁ>0�~��)1������� y:�+���+�$�PQF+ ��6� 9|t* Hu@�tWPW6H�q;w��mRP(�/t$�v۪m�-0&_kz)��Ϊ�G
�H��� |�� ��t�a��WL�������  �e���@&���	H�� t����HP�j�$PSЀ& �� ��F�%ϦrU�73�_^�#V���N����<)\O�U ��^ÃkOzktz|�y `"{z�s{u�t�qZk0 �q�qKkik�{~{ �r*�n,|L{Tr�{	�&-�n!" >#�y$�y%*'cL&N(,  Ƙ%l$0l$9l$���$�$r$�Il$N$�af$�qsSf0HdD�ye�E�yxX�`�ryY�~lffLMrRfZcC�k3�Ff�kAa٥ �d���u��<t`� �&� <tU<tE= w:�6�.���i�� �;	<3w� �6�qj��y�.*&��!<t<
t
�tH��O�Z3,	��R
E �`@� �#k�l�X2��]=I�à2��%D��2�%�`�j4��.�	w8 �wQPR��R��\C�
C�����.�?���.;t��>��WI��:Rè,V)�!Ij��MjA�S�[#����4k�'C���ziA	�	p�O��e�3% �3� �
ĈG
�t1��$~�G�u9� P{"��I�-�M��	�7q� �t���VW�wdQ3��d;�u;�`�r���r�	5�_��(+���΍��;��63�� �(	v'�A_^�3��tt���� �����AX	�� ���!�t���X(@�+Q���Q�0m�X&�TTO��;���u�c�t<o( m�u��uDB-+�MVP�5�w~�$����F&V� ��L���L�6� �@LJ���!����N�Z�x�Mt���B t!z�$`$@c6�6��� @����3�8�sS���"j~E-V=�|�ƒ��+�xġI���LX"��)�RBw9RJzv0X&��&�+O���͚� �.?��S��(Y� o$<
�u� ��z@�0�� 3��Q��)�ÜYW'���E�;�u�*kg��A\H�����w�@��PAu-����<��Yj�To���ov��v�����$��6�D�W� t	�9 uGN����2�UI;�v*�q�u}���4��GQ��ޞ��M�JF���'z�`D-PV�� ����f�T3���M���5$e$AI���^��<��@����p8�su���H�_��W��u�
f6�>	[0xg��ZE��t�W9$rBd �Yt��F�t����;���N�]��; �Fs�8 uC�����6��'�A�'��>�t}Y~�Ƀ~�n���FB8�s
z��
����u�w'@ȃ�J�� I�<HP!d
�D�H	�?���}'�u�ld��'	vW�ثx,~�.�ʻiD���IQS�*�
r$'c��������	!�K�x�'��$������n!� �N�� u1���t�i*��-���P� Bf��X
�_^�t���Js���nH��Ԍ�
�]$KST�\�3%����t��~��^��& 'r��&t	�����p/7�� u2�����uI�� �%�5Ҵ�o�Lp��("�
��l A8�����Lwa�b�'`��V�� b�t>��Y0;�s
��Tu�� �%���;���$�؉\#,+Ɨ�1�D�^��� s�< s,�����c���p���>� O�>�2�7�;>stB�p9v<���8�SPQ����'���LO9	x|�
7C�	Ga�� ��_��X�ё�T�r�NH&�O��$����w�	F�f�'\}�Qud���f&8?��N�I�b��p�;�rH�)� ��Gt#O�4�9m��uNO����tF���~'�=s��l^sR��$Z%��xsB��2�� �z_�D��Ɋ.��/�?��"�2q#,Nx�N�Ņ�C.��n��n��� MT�{��n���Ս^�N�V� >������ډ�u��~դ�X�P�k��;�"_f+� q��u�������C��`���M�6��d	ʸ�"����,�뙂.F'4�I:�*uuO�#X�	���n?1"O�� �!���tMQ&�u��@P=gH�"��5/1���x� 9*u���+�V�� )(��	N� ��V���!	�� �H;�s��q�댛�/|�����+���=� 47�$S>D�}~+��ǐ�M�`diD#�S;�s||��~K>�c*~"r�K}4��&�V�<S�b"e�/��;�~��?���k���_�S~ܦFr~���sT)��?*��tA�Ý��q�
�2?�ts&+�2�1��>�� �;���G�F8q��N����R)[[<r�k-�gH� _�������nn��u�9$�V�H�s��|��e5(41���OW�D�@������1��(.S�D����	u:;x�;��v��%� I;�|!9��>	w96v���;�s	��}V� F�q0�_P����[y�̥/�s
o��S�wd0��B"j�,uH��>� ��^��N��V�0coa�19w$�w<tO�u"y;�t�G�
x��WR\�:G�>� 
�u�7��	�;6~qN!W�/+�0#_��>���+� �tt�.����?���=�
�
�&�n��W,���{�D��z²^�#YE)6	�s!T�
�e��#����L�Q���+Cxw%�P�"t3�~���y�����#N'���Q�VՊd6 +lV�����|^��8c��������ŕ����Hq(�����z�p#����)~E�39�f7��]p��;(�s���fKO�4(������W�
q0���VRmp��X��z���zd�� BQ��u�Q%s0S���

����(&�^�ot��Vz6&M�J�P�����m��`! �/ ���)H 7O��K+�L�!�c�u��vG��MW����(��&������R�EɿE�P^��K���C�&� \`�t88�� �>�
��6�P�*���A�F��'n �v0��F��&V�\�rT�a�},��[�-R�#)w�\y��� ���"ȁ��V�M�t�6?M�:er;.H+�ɺ�3��QQ�	PQR����.�V���t��W��^�WD�WNF�x:'��J<u7M��QJ�&#-�J]PH�*+N�.�����Px�;�s�D?
z� ��9wH�� \7K��"�u�%.dx���ٍԶ����q!���˓03��t��)9	AN�>?�"�;rq�Q�������sЭ��DЄ$>;�[�zQ^�P�X��h���� �&���|�YfIDs `�s3����+�;�x����+�HG��K �O;�s��\`/©�+z�
�'wC$�_��$n5;�8�b�
�HH�;�v$;���rr�M$n�G����O�X?�w*�!7*>�vb�xN�ƣ5�"#�vQ��p @�������Qt��|IKp�!��$j��iI���.����T"P�
�B�uas��T9E���98 �uWH�*�Kt�W�r �<�����+%@��.^$o$�Z�Q ������1����+��4�ls���V&|K@ء�N�� �	Sq�oU	HE3t�V5��妬X'>��_��'1�Rb|w�!c��Ñ��
Ec��^��N��V�n5�"�<��ut�b&���"����s����#B)7�XkR��Y��Am��� \��R� �+� ��܂ � /� �t����t�+^v1��+Bb��$��9Nw��N��I�!PjV�+	��x�Gأ&]���ʒgWG�����-@*���<x�F�/�*P����fOuЋĸ�ķ�wt(%���
�ZQ��3���E���	Ϸ� r�>s��t�f�>�S3�u�.� ���`����u�9��,	 � 	���65� ��GSV�� ���[YSW�H�Q�-u�<��6X#�X��X��2��D2����fH]�X\����6��- @�&�&�F��-�=�
s0 ب �yÊ��~�F�^�N�GG��0�8�� ��GQ��C
�  S7� "��% ��H2�!ãPq)>��pB����mW�9��@ 9@���L��� �(�w��8 ^0�%��˫�20D��� ����t�u�BDW;�D��96�u�D���&�>*n���a��@�}9uu�E�.o>�Ժ^_�~X�f �E�Ʃ�D*D�f�E			� � t
�m�m��t�M�5

Ql�
;F�Af�			VT�p3%;%� �n�?Z+S�&(�	V0 ~�Y�-�T�D�r6T
��3{	aa�as3-		�	Khw�Y���������p,���`MF�8s���}.�.�%.��|	6��uި;��,/����
��@����Q��+
�� �xG��u
�r�d C��F*�P�J�R����3�	��8�v=3�v5
-�����Μ�Ν.�JPL�P��
U�@e� �'p�k�ԧ`/��5���̉��*9�Dru,���W��T'*�H���G��G�D	Դ��Vj UPV��/�.^G��鰟L*�D	��A'w�����&�� ���N*��s��L
��Q�*�F<�KE�
�I
Ч�TL/�
��LLP��Q�	�9����t�O�PCT�|^e!�5$<$5�,��u,0u96�uq�P�@t�� �N���XcP���2�~���41�5PP2�:Ý�B%�п�Y��� ��2��#�h�9�_8�=9����y?�G�� �Ts�hCV���p�Ї�BOZ��8��8mML$�w����9�
��TMH
~�Ǆ^\�E�A�n#=V='o/��+���V�A�P\���4,B.����w������ �u��.D!H�{LPT0 X!��-������@6��sFG��L�؎��N;�r!T!���w$rF_�)`��/��Ŕ�72����;�uQ;r4�4/��/�C�^E^�>2�	���U��O�_M7(URIXu���D  ��3�����A�ً�� �3ɊD�&:E�OrI��I���9W�A1/@��_��+F� �+^���ޚ
 KÃ� �N0!�����(�.""�j�u3���B�� PP�es�DP�	�.�WW�^]���{ �uu� ��@�@ ������.+ ���!�  r8u>M�/�� v �� �V�?���ڋ�7�,+0tN������O� ŋ�:3Ki�99��t�>C���&�]5�0A1�0�� �߀�A��++��:�%UB�XN8 	%� ��D:\�t�0`$,@:,t�дG-,i�V��]w6�|.u��"���.��xX+��t�;9��s���x�q3�b���� :�6h��P�a�3�:�uAZWh��z`�����)�� ��<.t�%G��?t:���X�II���� u�����E^�� ����@	������VX<�8�< t�����qtn�r%\� u�?..��RĀ��j�/naV�z!`
[3v�F�5j4=�0��~==` }i�H�w���4P�7Q4IeL�,�,p�? =�3=R�\��&4 �$<t��`�F
u��t�9+t �DӃR9Ku��g��g�g���������������
� ==%r���=&v.='`�ax�=(%�p�/�z�x��L��� ��B��OS�7�4�"�*G�==�3�
=�>�h<��~�#�9D �V���K�Z�m��p���{ :a� ��{���7���9>u��':�>�- �y���
�]뽴�����~
�A��S�U*-�-��Ysmn$?<4d�=% �FW'����-͋�T2PC�HDP�p/ 	��i���
rS��g8§=������f�� ������=D\=�&X�= K�hM"H=����Z�
�*D�\w6jv�> ��� �e!V�d!P��.�[
j!��V8��"JrP����t��p����$��t���^��q�*���G���i�`�5,�F�*�;w	xD�F�#���+
@���� �$���  ��> � ��D$���/����Nd }W�^�� �O�|WIS<E�H�aBuk�>#��u��d���;�tT`��S@�XSI�"0� 8= u��	?c�_� U.I	�2 HH��KH�H �Od�R3��AV��<G�ң㈺6H�i��>j[^��a�~
d8>|� u��Mp�u�E�\���l+t�q-{�r�%y]NE��M>ˤp8 �b|��׮D�:I�V��)@󐓒%/�|�� t9�>�-27���E
5�tD=���[P��]t�Z% @W�c�N��;�N�����t�ە	�b\�	[2������} ��Wڿ2u�,9�D+��V�9��aU�d���t�#���gj�V4]VV��FΞtT��DW�Hu���	�k��=H=���v['q �F��f+8F
v��&�^2��R�����mh�FN� (F�J+VQR��0 6�>�������t���u	�w�		t ������ZY^6'h+�N����]tj[��kk�������o+�.�}��sF�:�QW�_Y�>*X���6�>Yb
�6�6�|d+8!$��`'�u�<!O��PNn 4&���1�
W��F������D4WG�O�;�t
ͤ�W�% �D$��P6���&%�<�dYs�KJ
u
�\����O �F�%	S�5��$H7<O�V��ƛ븈�=/�=\u9c�E�G�@ u�Dt%�Dxoy3Е�8��F�M�:V�a�h���Ѥ/
���~��&� ���5�J��p�G�=*�vE.�=:��=?�\�/$��.B=~ЊD����<��BU��]ݦ��buTy�"#8���p!�U�;rӡ=
��B[��FG�wժ��]GZR^��A�I3�V�P��Дo�q ��� u3�� �]�\F/C�-+:�a�)Y��� \.r>�I���u���t�.u���H.�D.+�vǽ ��G�}�[t@0*�=-uq�F3:��t�!�G]u��w� yqKp֥�"�4��*�+��`����;v���7\�F��sw%tOh�O�.\�:OI������n�+�����"N�"�\�u���b!����
��/1��<:u�� D��q�*t�x�?t� tH1�F�Ʀ�N�9`t�O�|�`
F	����\�</u��.t���1�!N
p��=�A��u�+��N�+��E`uVW��>�`�� *�8�>l���D�D-�D���0�=�dFq
F=~�^�p��;u�B m�L�u ��}~uG��6��*ɀI�*�ȉL��%�����YL �ŵd_P�]��tt���`�, ���v��0��.��$�FNsht�)��?���?���U��mW�]#�z��_�����Fp�(�(��=� ���$�WP(%v�K��p)������\�tb d�tw�G.^�*�I�RVC��(��$C^&=}�ħM	t�R�j��5L:bHHI��=�����:N�vƑ�*���$�v�@m���䦅z��t!N��^@G�#�P�	݄�G=�u8��}��-&�t�k���^[�������?H� t�S�����PБ�z=�L��uL�܀������������pl����kb�@�|j�[� .8�鑮��r!q�  ��#>���c{�����D�u<l��E��*tҫ$P0.}�@�֋�$:
̋&��/ )'���j�F����1��u��6��)��{,�RP���5o���F�u 7XTLXR/y�HA�!C�7�~�.u��DeB1~�&1'F
u0dBq��{$;��˓[Gs�z��ou��� $B ������\>��K85T�"�"�*"ʽ#�΁#"����F�A�T9��Rw��>S�l����Z~�,#�N~  +++<<  �89:;<=>?  �� T&&���Q P��t %�I;�PMd$+$R%@2��64��6n�HL+*M6�H��2$0.�>�p�	�F`�8gt� ��_��G�E
q�.R:F�rU�  �H �E
@t�.F<Htp+u�����S�0�[2�5���6�G
|t ؊��&�&��@ "1&��M �ub��Hu�uQ���+ u��S2������Y%2u2% t,�3���!��	�
���`��L��  1�  �p��	�E&Q�"^���� ���- �	`t� �@%���` �~�d$��}L'�E828�`H�E�4�M
Vp�׍}��ؾP ����.��'"pa���@+��@�$�f{`���3�t�  �&u��e�6 �t�}r� U�0�3�o]�U ��M�=rw�:/6�a���9� �:Tw�����`w#rP����fCXCt��q �9�EJ9_'�DU3� ���7�� �1J	1��Hc[VW*���U9��*�� gF\  t�}$�; � �X��B��~�< :<t<@t<�[< )s�Z�q�D�N9&��G����
��a6��}+u�ȴqb���1 u+��2KC� ��� �#2����.���E "F ��צ� u�̋��]�-��Q�����%M
��=�+0�9 S-#
�x�MO\T]">�P[�_l&�f����R}R`R�>7f��#$�Q t��c ���e ��� ,�!�:u 4��u©fB:U�K��
E�%�:�6q�	-P-�� &�&f�0$,t������&�6��ãS�3��X2�P�}����E\CPop4H*�-\��<t<���B�<�����;�~ 0
���� ���r��w��� �" r�{ ��� 2��mO� ����d t� �2�S~FF����' �6�G � �f��P�7� 
��B@� r4�6
� y�}U�Ө�ً�3����'n^t�`��e%������� �W� �a���v�
� �� ���M 3��_,7e�kP�L� Y
�

0
�����C9 N����@ �}����n5���LM��M�������r"3ú�??@�� B������r<t��<�����7�X�r5�<�� ��K��i���~��`[ t
��	湑[6q(3�0���@$���o�;@ ����Ўظ�QeQ e���$\$�^9� 8E
htz� �? Ht�& �%�I��V�{PSw�.�7�9 ��.��d+�� 3��_����5��`�!S�%c	�VZX��
�t��f*�~t.�:LZM��
�u.��?\���P���tX�0�S���; [�/>K"���qCO��Q

O��;w$Y ��� 2������_͢x+�K���W�N�1��.:Du.�Sp�|t
 �dt	��B�ߺ������V˜�!F� \ ���r3��� ��������YjU޹ �:P_�4f3T^]dc@��� ��@�0p|�Tt�U�.�`�T�U��eG�5T<�7
�3���`D�E�uY_���$�}� �&�� ��S [��ÊE
�a e�� �U� <u"-	'~tY\~tT5'<t�t��pnC�� w ,3�t;�$0Ѐ82� u0$��-�f
t�n��nA��	th�
�u��Ћ< u�����E���Ct\#) �#%<t!�.�RK ��B�� @�f�������Z2���;;
�ʸX_ GH6�3D�n�ʀA�� (���|t8S� tPA�Xu'�� �����u�X� �	���u ��[�e]�2���&�u�@��Jy�.�@�t(�͵�8P��&e��xL��ސK^�D !�v�V
 �h�  �M`�r�U=	o�2�6�:�X�v��ψV��6e ��������2�X��O�RPQ�j ��X:)?�+�E,RG
/B;�M�c� �����=:]s3�N�*��n��ߺ �%��0�5 �"2���ܫ�����������t����4�2��fS�pCZJ�
#`��� ��U
�ZÂT�f�H������uT� a��X��� ��g(�!��߬��Q���`���^�	4�l�LW_�^�&t�s#�D�d�povT߈E�8E?�I���	  �+=$&!m%'k  #("-.ghimdefkabc  `nQWERTYU  IOPAS D!F"G  #H$J%K&L,Z-X.C/V `0B1N2M�0�z�{�	  \[]';(')`+\3,4� .5/�-�=s%t'u#  v"w$�!�z�{�&��( �-�.�$�&�!�%� '�#�(�"�-��z���{�z�?r
�t �W��t�ʥ
�9�!�Ǹ� ��U;�tKP�`  ���R�Z ;�t�RP3�#xNT�XZ&�	3��5t� ���Ӄ���  ��u� ���
M�E��PR2�Q��Q�W�PSOGZX��q ��$~��$t2�c��2 M���G�v�_��2QQ��Y;�u ���}k ~�En�p��Mk���tn��C���_�O�lLv�����  ���?�\;\�Xv7�W�Y����2 ً��AA��;�R�q�0�1�� 4�)o�a�$��~�2L�(�@��K `r� D������`�UP��� �7�6� T^mY�G��q6�d��B���E0�@� �E����U�#��G��M˻n��5KMF���  ����O�g�N�
�����:i Ekx������c�s	�ź=�� ��Ƹ�6�&�Ef0b"` �n&���l�E��:h$_ �V����d ���3�uC� ���U�%��!�,6
��#	�		��	�}rK.�����롸 0`�r��=r0 ���r)
�u%�G�0�)5.�3 �.��� >�Mr�RPS�!��[ �߉�GX�%Z%Ã(�v�ٔ���0��G	�qt� '��_���V V+3����Uf2�ufu	�%���2��W��r�^�3ۮU�x ��u��SQ�eh�� ͜�]t"�>>�	_�Y[ÇO���)�^J>��.�5��<q �:*�xX��*�R+ Yu�`�>�@�e  �Ee�t
�Ef&�e� �-i>\�Y�C��D� gZh������ <�6�d<�td$ 
�y:Eju9��i�A on�| ~'Tj~��S%�`|0�L�Mkm p�<9u�Mf ��8�ef�� ��o<8tk<`tgf�a�'<Lu uX׃������
�����'�;t9S  �؊Ȁ������2` ���tt���f'�
� n�.�[t&�S؈ee�=ΐ�D8� _2 � Ü�L�	���� ���V���u0�\�g��J�p�u�Ef�ЇEr3��������ى*��^�z8��u�8HWP.���p���
 �|V�5�DEk�}^X_�PP�6-VRQSP.�.s u;�1�tH(�v�s?":�0Ntg�܍6�gX[YZ^�)P��-�y��u�lt���fo�d�9u�qI
�����XP@����@Y�  �6�'�6'�.�6�����_	�.���&:��u�_�
��2���#�ȉV�  3ۉ^�3�
�u�M� p����u��t	 �u�N�����,�F�9��(
�t$����,d�=�+t-t t��� ���jM7��k�!Nt�mJu��K(��t ��at�t~s�	���~  H������<Ar<< ZwY��<ar<zwD�, �<rܞw@��.B�� GɁ�u�-k ��u
2ɳ6��a cGrvTsq��.�n�1�s� �N��u0� �B���=+�~Lu!i�]��ru�'!q{��W>3pMASu������0@ʔ�9w��Kt�8�x��OJ�c�3� ��p�;:�rR>Dv?�x�T� D]v1C4�^�3 �gv 3��h�#@nqv�x  �w�1���Ċ�	V  ��T��]b���uK����t�N��<���@���. 3�����������kFE`>�.�����#��� <��
�t��S2�E.�˟R�c�P�3ۡ�v�$M���rÒ��>dz Iu�� �E\ĹL鹬�#��`�C���BX�a���a�< Q�0&-Y��$��#�l��gˉ�=�V�q."��!� d4c�  ��> �!u��` �8� ,,6Fjhpi  qjrksltmunvowpxq  yj	x1y2z3{4|5}6~p78�9[�  �	��&�%�(�m�k� n�$�z�{�'�^�}!*��,�.� w+�-�'�/�;` O2�W^  p_q`rasbtcudvewf�-xg� ō	�&�g�h�d�(�  b�`�.�-�n�z�{�0�  1�3�4�5�7�8�9���f^-
W
�@p�=�;�'�,�.�/v	xI!J$  O#Q"TpUqVrWsXtYu  Zv[w\x]y�&�(�%�' ��`�n�z�{��hV��0�.�6 H7j;p<q=r>s?t@ 0uAvBwCxDyG$H&bK%M'dP(fR-S.�͘z�{RN�@*SWW�Vy�(��y�����(yVEy8y-��y�Ly���'y�a yG�P+EP���P�(�P�Q@P��� �d�IzP���)�P�ɥ Po� B��wP(�pPT��2<BG2,�232B�.2@��2���2M��2��H2~��2r:�r2�ߪ	�5�Z2,J�2�+2� +t2� Wc2\�2
2��2+�#�xS��R�	�K�:rK�}#YGю7�#�(#W�S��G�O�[2.��!d_�ifBt&} f/t7t�˗�^��v���uK��O	WuK��	�tY3,����971OH$I3QI9I2I5L5���
+o#U
R�
-Sd�h�f��q4�7���� R ��u�+�k�+T
S�uHq�-�mu� iV�z����|������� ���F�1���T ��������t%��jt<Ok��m��n�<�`��� fu]�V�A�A:�rr�Zv/�a�zv$�v�0^Ȱ0W@ǯr�`
>*�*��2ۊa��.Vu�Fn�_PZ����L/F����� +���<��:��^&��u���̸Ì�6�8�;ʸ\��U>@��<t�@��ǅH" ���~�x"w[�^�8��7�F�2�b�B���CK<��Su���?)�F��V����d��č�t�
n
�5d3*���P��~���PP:�P�B�PWA}�� �v$��3�WV�F�3��H�U�Fߚ)�S�h�:3��N��B~��^�������F" u�Ft��7��LN�oV��� e+��j3�GA�sX���MA��Az��6d,��"��^6X&��V���GW��V��=q%'�� R�v��6�|鉃	�`�]� �?	u��f� �e�b� �-��# �&���v�B�B��X��ua�2&�GoWq��z"�9*5��)���C;�9��$��a
#m�����[�I�)�+��������>>u�$��G3r�> ��!�0x����7 ��!��  �H^&;����P���f)zV3/�³��8F"��:ڥ�(C�������e��|�b�9u�r4(�
��@����v����r��� f��N�y�#��#��P��~����2,���B}�)
�<Ȑ d���Г��d��Ѹ!��D�]�h,�^�����D���FN!j��F
bF'�u"��rB �+ҋ�V@�lP�
�7�4�+�V�;2�g�<S�`�Nt�yH�H�u%"%���'� p>
&�l򝍛��T����P.�G1%v f��k�F������8	�#d�&9G7v�"�c��#�1a�H�G;)��*+ɋ��}<%�p�:#�/�w+)����S�@����ВI�t=0�e'�	)"R��W��T��~�Sr'��ҽ�f�V��gt�����A��F���F��͐�VeH=q���� �����@m�FN,�
lj
&� �~�j��7e�"�!ʀ}�G��ǻN�z�i���8V�)�QI���q8g�F��3�9o���@H�c�n��F�����~� t�a��^��v&�8>u��L�1v졇l���P�Gm��EB'ƴl�.`�t�64�����5~ƄdF�d&%����|� d���]���=����:��=''��tdb���9F�u\_�5�
�P)��5
pE.,,PQg��:{��xa�S����=h���w?^D��S�yu ���&�Gs�����
 �LCA��xn�,��K�Q �<qI��"x<����!�=�	(z�  �z� �F�t�����0��-����M���Q�O����uM)�)N;�&�͔S�Su)m�+�;.w�zr;�w
��D���+�	�j2��1uI�a~C�#���5�t5��/h�{��x����s�����R�gb���YԎ">�ƛ*�� F����~� t�����	���&,��A�! ���P68��A�E��� ���� ��939��@�3��b4�9F�r��_u�c߄��?��.o�Ij���� <��F�t+��t
Rtj��|�����y_�r�r�CH�O���*�ɉP ��	����V�G�XF���1�� �ρ�ဋ�%"�FI"k���B�`�G�x�B�$��:����	��	�}*$�$�Rى.�|,~��t��ދA+�r5���� c�^L�YJ�CRt� '?����N�&�;�Ӡ2�����R�V�qYZ(M?�2�Lt��N8���
O �U"H�ldA���Jv��Q�����BH�tV=!�!J�H�B�r�۹Q*~W(�
r�V28wL�tf�EV(���Պ�B�V�K���D��lՂ����0݆R�V F��^�~�&�U��8 KE�~+�ML��>�tX�	�NqQ�}"QCM��7	���+�I@�0��~��:	-~�O�%�~�$t�:�ɘ�P�r��G��+��9�=�!��7��X?n!	!Y�
9�WV���~�̅N�F�۝�IJ��<�IKK!�*�����G��A�S�'Ha]��l
j��"��Z����rRU�	g#5v8��3m���7�KN�NjR���[�v�-�H���@-'�e���� ?�	�Wl��g�!�����ڹ]�x&o$�X�t�E$6�2:�VH�� H�����8���⋃��(t	��p�Y��`��Ƃ�� ���-����������>�����l���>�uY�
t�� MuJA��;�u@9#i�,u:T$p ��ؑ㶏1	{.�_�+t��]��;+��J����o��y��~��uY;qM�t����@ �*���s, ��+�h�Đ�^&�7�#Naፂ��B�M+	�T�1��	��	��L�gѷ���~��J������d�].ܺ �� ��Gt+n��*�H;Fvn�2�
mf�n�N�tJ0u&0�?u��~"-	l(@�+�1��&O#EYx��0�Z��̾�ǿ}�Bi�=>��j��Q�:fV����Xb�\��f3�HH!h6���|6"��Wn)�!������4
و8�n.t��u�/��G;Z4��&��-9|�W8o�
+(���V�ĺ��5�F���B��F��F)X�Be��p���F �-�/X&�x�"ۊG<wr���O��Ws��;�0����o���ԥ��&���昞K�� �H�\�{�&��D�!���tڋ���y8̣���* ��"#�#��%�ny?�� HF�n�i�x��h �w�9	sCt H�}�����;�s� ��t*��v�z����8FG� ����F�H�� V�8S	�h�P`� =�u�
� W�*�u���9v�v%��ɹ4�V
���:�u�|���7$��}���~=��	�1��|���8�  �zFo�� 
�VW�v�  ��� ,<
v�~������y� �| [�.��(�e`> �CQ� �Q���S <p/�>�Y��+��� �w��2����Qm�ǰ�����Nu�0� �-�����^G Y��&� G��X3��_ ��F��t/�t��� ��^���&�5G��u�V��r�
Ö�0 �y�%����ZT��P@PR� �jq&8%ntg}
�N� %t��u.w*� `��&�<Zw<Ar 0�`%G��=�� :�u�`(��F�$t"H� @|N&�}�  �u@��� t	tA*tH��߼�] �����I�EJ_�p	}8��n���˲�4��^5��@H:�u�N�ږL!�fW:=!�_[XY3��R����[Z@�uAuDIH�����X,a<w�, am^x �� S2�7CC����+���no,:' 9&9Ow&+A& '_���� 0���t*�؀� ��&,C �g:�t������C@�/��
u� #:�Ht�������	�g+�-���k�e�K	+�8D��t�  7
l(� 
 � l�31�03	�b H@  '= ��K3R38 ??0�~HelpP:��nt�H 0:~U p̀f �/� a�c�� r)����{�kW^`^W]come to�hMS-DOS Edih-r  QBasic Copyrig`ht (C)rosofrpatio�n, 1987-92. A�ll 0sese�rvedPE'ntbee�Suiva1G�uide&SC��$clea-hix�#og box����C  �Z>�
$	u2�#�d �C$-
vm@�0
�8��� @ /n�g420v�Fi� � ~Name: ~s��Dirs/D�v	`�*�7���z�rݣ#���'�L �Dr�	��"��9 �����	��"S	0�a�h\ tꌔg�q�{��e	�����
�^ �Ȝ�y~S  vected Text Onl7�y����Progra� ur Win�dow omp54 Do|	cum�5��;H�8X��D|1v@�2�~��{ �   !�)��	�	~(@] 	����*	����@�i��%�c�topicCz[$#�on
 %LPT1 
n�| `9tup.� 8Q (�``��X  6�H�
�Ml�j���fQ.�
��A�� T *'���Us�ap�c��n��T��~12��3�OM��C~2�BLI	I&e��Q�@����o '��(t�' �P��Fh�ߒ8�Ja!��<6�PZal,FBKNN/���M ��UN�Pr,D&	;	^ALmChoos��V i�mu*Pe� ��n ~Act���ee�:|AU<]���[T�eQ�8�!DL�&@���iz��
яVR�\ѯr�W��-0�N R 1
�SQj� ,+���vJ8	ԃ 2E&�1�2� ��o )	HY NColor1QC1. 234�Feground�BackDisp �lay Op";?7S9_#DTab '*SIsL�D.g�2y:�o* `"�����KHELP�*:�`f��6
+D-�`z)Mi�\N�|�y$��k �t 0$�(/q�iF� W�8hat�Cng�sTM `ch Upper/Low8�casc*oH�Word 7F:2~Vif��AB=t
;�%��,'��*��D�D$Ɛ@S %��D"�d�G )"��ξ
��0}5Q%N���0ސ�]��@@& R5(mf�G����kipL��HJ�\ ��<<FMSG>> �R60�#
- stS �Fov�fl� *�2�!X po{�no�Tded''36'|]rFv�'e by Z �!8!9ea6ughopo#��f� arg�Tws,	,9� ,Zron��/..1��ill{(��n���useR�&&3z�&f%�g%4%N��tA-BREAK��ru)J��'5'!�exp��Irup���.n-ti�o��N�q� �#'�Z�=	L	 ;C_ �FILE_INFO0� �3F�� .C �psqy0*4*�{:*�"��WW *d�.sc���4�O�b��c�rc
 `3IJ�C ^Lc;��T3#"#V3�s�Fc@� 
�PO�?o*1찖�D�P�+�LE�q��*j-���r�Rr%�T���rˀZ��t2�q�r22��L�1��New�pen�yKSa��� AsŔo
Ex�Z�L"~ �B���N  ��	���c���t�� Q �{U0@p@Cut	Shift+!�M�3/	Ctrl+I���Pas�BC�	�(ʘUB �FUNCTION�C ! L@��Z�{��Yx .� A �>����p )	F28�8pl#O�p�p S���4dL��?>��|R��/�Rep͋�2L� SX53���$.2/&�w:�'N�t*`ar6F5^VsW�>nueV��),*ɼ>�+���<�� 8�ocedu��A10�Tr�O	�gTogg��Bak�U!9 �[�f̈́sRe�N򗚗B.m ���n1�T�u7�x�Uq �:�<l��%  ��&eQP[hSy g`ax Check��� =:b�5>pn	�es^( |RT��x:� �a	�Ind���2� xs�`lY��$AbouB�^F�FC�|��E a4� ��H�G�Get	�\�ed Key	�La�F��",�G�<:Ho!�wpR�Y�J�I�� f0�$9���Vi��8�ich2Pun�ebug I�F�p, D��"<�H	� ��  i�� hm  ��� �r8J~40�0F7�P0�@	t�@@X�0P~���d��6���0 ��@Hc� � ?��" �M�P
�)�Z�HV��D �+Y �=
-Z 1�cV\- �& p	^ ru��J�K�GC	��E N	_ BN�Lq�XDs! tn5+�)��[hvS wz�0x9 y1�\) x�����H�S���l�@L�RUN-�OC�i�\�B��� MUr tl������O..*.TXT ��\����y{m�Rqb�.i�ni;09.-A� Z-azB������� �����������
�& X� 3�  �O1��3���ƴ,�  !2�R3��Ʋ����&@��
X2��
������2���n
K� ��>u�۶�(a�Eu͢����< m�/�g�#"F��0����6���Ґ���
0�'Ot$2��O��2��+��O�sa���6PP�2�Σ �[P��	3ۊ`����a��-��X?:uu:wd~Ê�*X6�BT�X��@=x  �t�����]˫��߀������� `��������߻����ߵ�������*߳���߲�00���������� ���������!�����������������?���#Nh7�@�>	m.xeQ�
a�� � Pd�0�.$Q�gR�P Q�^!�b!��Fm�xI�a
 !(INCLUDE��h�.Hpxpp�[� fpGOp0p?x/?
�1* pvNt�c�B01f4 !�o�6p<�
����Ow��/ F(r� 	�=	0�ayu ptc_b^q wo`p3�xvn@

�7DKBK �eigfjhkl_S�Y��54� �����-��C� '0��DBF r]STA TICDYNAM��\D���"+ R
�d��NMp�ALLOCP� J�R"�,���E̬�Ult�����3�F�
		X"4	6	ABSO�TڨE�n	�=E�� T��@�8�6�z�z
� ^�,}�`W_QB��C=PATHLIB�%q~}�D��ʾʐU 0MȾU�U�UL\�
]� iMBAS .E�XEL�^�nJej�Wqt�P�Z �&�O"aW��' �W�xO� C�3� ��;(@Ȍ �d�y�M�n*~( ��w � 3��Tj���������| �d2},�o��}"�$�6G��nF֧1�"���Fd$��i�Ce322&�1#NANK�YDc@@f$�7y�AC���>5�h �!����?��pr %��ܧ׹�P�fq�@� 
�6C����?!#�p�Xt�ʄH iI*H�IoIlI4�#HM[H��v
�V9 �VIIlH�I���I�� [��|�9�gU�HFVH�I��s�?MO�ଁ��'�J3�&*RJcos�� JFta�)0�,-O00�H 4J0IaZa�	R� �0^H�@a
 �J]K��GH �0�K� 2 �J�K��*HfK}62wK �[H� 	�.���:�I�{�$����J^>r�*�JQ*p��{�
�L���I�j����g�ym,s�;������2�+�!��!ɠ!x���"�r�"<C� J�!(C� U�"e� r�"^e�!�!W��!q 4r%a!vu�Md�l��M�'�/A.)�I�8 8�H" �J�s2 37�:�WX *�OH�a5�hU�l
!��
�j��ڿ���  ĳ�ôɻȼ�ͺ� x�� �	&-� -	�8O� <c���{5�[�=bij�c�����K8k=T ?()} X�[]-�* ���  Ԉ҅��뇀�������  ����������ӡ֍ތ  ׋آ�������Ǧ A�I����O��Y]��O^Canc�� Y��aNo#t�try��{�6\� `�NYR��AH(� �1��#*=��ov��[..] [- -]P������g��!N 2f< �& � �,b�<�8X"��|o�^)��+�.�3�a��k�`yF�6��c����Új�1�����l�c8���\��3��_�ϼ�L��-�y(�P����"�gl� ~ #����?�˖@� ��@�5?5��<��� �1�B	{B4 � ����Ҟr�?���A�V�>\ 8��C Þ&  s�K"+,:;<=>[]|  ?@ABCDHKMP�?R:EF8*6&#{��C�����<DI\R> sSPEC|=\	MAND.��C�	�ep
	_ ������<p�<�$8Q�9X  � MD�?RB�� 3�� �Fo  ��� ��O����P� �4 PˌÌ�H�����7�S�G!��H������H�+�s*+ҀT����ڋ��*���¬  ��N���F��$�<�u����<�umm�0gt��2��x`q�3�)����c i���t&�� ��� �t�� ��[@������an��>�6�t�3�-������� �����.�/�@��` �ʨ��!��Ln�PM��f�-l  ������ã�r�-�  ��¸¯¦�W�6  �-�������y�\��  ĞţūŻ�������K  �sƒƦ����^ǚǧ  ��C�XȤ��������  ������&�̛̠ͩ  �z�r�f�Z�N�����  ��˨ˁ��ʷʒ�X�  ώ���͒�p��л��  ѡ����� �E�M�q��  �ԀԎ������?�R  զ������<�E�Q֟  ֲ֭������2�D  �W�~ת�Oقْٰٞ  ������.�pژڪڴ  �ە���$�(�����  ����ݼݠ݋�~�m�V  �Q�>�6�&������  ��ܾܲܩܑ܀�m�h �U��{�r�A�9�  �����������s�  b�+�����������  �߯߈�������3�  ��[�E����
��  ���y�p�P��D�	�  �������������  �����������~�  u��E�O�����  r���n����\���  "�����Q�!���  ����������5�p���  ������)�E������� `��o���>�[���  ���y�b�:�-�����  ���[�%����������  ���(�#�q��������  �~�Y���������"�  "�"##-#2#D#s#�  #�#�#�#�#�#G$�$'  %�%�&�&R' )/~1�  34�45�67�7U;�  ;�?�?�?�?�?>@O@v  @�@A/C�Zz[x\�\�  ]�]�]�^�_�_�d�b"  b�j�jBmm�m�m�m  n�no5ooq�rss0  sFs�s�s�s,tCtVtc  t�t�t�t�t�t�uWv�  v�v�vCw�x�xFyZye  y�y5zDz�z�z�z�z�  z�z�z�z{{%{2{>0 {I{_{�{�{�{�{  �{�{�{�{!|E|a|i|  �|�|�|�|�|�}�}~�~�~T~q  ~z~�~�~�~L���  E�À̀���}��  �˂�s�i������	  �k�|�����_�}����  ����䋡�
�M����  ���ۏ����  �u�����#�.������  ���f������+  �ѕ�������.����  �{�[�f����Y����  ��k�|������8��  �����:�O�q�y��  ����`�i�|���̠  �����e���T�Z����  �ʨ\�����"�?�]�u �/�J�\�Q���  c���ʯ�'���	�  ,�����ʲ߲�S�t�  ?�]�����8�N�q�  w���ܵ��/�Ƕ�  D���¹5�D�K�����  ��Ļ@��������)�  /�=�W�g��H�ؾ�  ���B�M�������  ���mv�U3  p5 �6������;!\� � O  T����  o],�Z
 �����=��� �N7'  �_��_W  ��v�{c3  �
�
�
�
�
�  
�
o
V
$
�	�	�	� 	,	�"�&gu  ����`S�� �ՆvP���  V6�P"��  xQA%��P@  ����sG1  ����`T  ������  ����_'�  �����]#�  �!*##�"�"�"l  "Y"8"#"�!�&O&&
  &�%�$G$?$$�#�#^  #*�)�(�(�(�(�(@  (�'�'/''j-Y-�,�  +�+�+�+�*�*.�/  1�12}2�2�2�2�2  3�334A4M4Z4�4�5�  5�67�7�7n8�8�8�  8�8�89<:�:�:8;�  ;�;�;�;<;<<�<�  <=S=]=�=�=�>o?�  ?�?8@h@�@kA�A�A D�D�G�G�ETL�J  �LP3P:P�P�P�P�P  �P$Q5QHQmQ�Q�Q�Q  /R�R�RuS�S�S�L�M  �M�N�N�N�N�N�N�N  �N�T�T�TUCU�U�U  �U�U VVSV^V{V�V  �VBOGOTOiOzO�O�O  �OeW�W�We\o\�\�\  �\�f�f�f�f�f	gg  gXg�g�g�g�g�g�g  $h�hbiXj�jl4lCl  ^lel.nfn�o�o�or  rnrvrsssss  As�uv(x=|�~�~������  ���>�F������Ԉ퉈��^) L7�������  ������a�m������  ������"�)�j�s��  ��;�F���˹?����  ����*�߼����E�  Ԩ���g����r���@  ۧ����8�����Z  ���� �%�%�%�%&4  &P&W&]&�&�������  �G���:��^�v����  ��#��Ȩ��x�y�y�  |~M~R~���0�H��  ��y�ʕZ��������  �a�q�����+�K�t��  ���ޢ'�~��������  ���<�v������  �����ǥҥ%������  ����!�h�{+>�3}  3�3�3�4(575@5F5P  5r5�5�5�5�5�5�5  6$656X6�67E7T7�  7�7�7�7�7�7�7�7�  7�7�7b8j8�8�8�8�  8�9�:�:<�=�JSK�  L�L�M�M<NoN8O�O�  O�P�Q�Q�R�T�TyU  Y�]�]j^�^�^_!_,  _2_A_U`i`�`b�b�  b�bcSc���  !>Gdz��� ��������
S ��u�  �O���6;s  ���c�cIk�����  
ҧ����&�7�E�R�  X�g�l�q�y��8��  ��V���=�����6� ��������W����  ���ӾӢӄ�h�L�m  ��j�_�Eʴ˜˄�l  �T�<���|�P�z�X�>  ������n�� �$��  ��� ������  �� �$�(�,�0�4�8  �d�<�@�D�H�L�P�T  �X�\�`��������  �� �����  3P&8�	�\ n��\iA _��@������  ���t�R��~�  �<�����w �W9_��� (�pJ;��  ���?�A��  �OE����"�  "�"w"�!�!�!v!X!@  !!!�  �$Q$2$�  #�#�#�#�#�'�'�&�  &r&9%(%�+d+�*f*  **�)�)�(�(�/�.�  .�.�.�.�-�-�-�,�  2\2K2�1R1*1�5�5�  4�4�4�3'777�6�  6s6g6;�:�:`:A:*  :�9;9�8t8K8>8X>�  =�=�=I=0=�<�<V<G  <=<�;4;tB�A�A�AW  AA	AjE�D�D{D,D 0DaC�B�B�InIfI  �G�G�F�F�FtMMM  L�KGKK�J�J�J�O  [NSN6N	N�M�O�O�O  �Q�Q�QR�USVlVtW  �W�W�WX'X7X�X�X  �XgZvZ�Z�Z�Z0\d\  �\�\[]�]�]P^�^�^  �^
_�_�_`` a�a  �a'c:c^c�c�c�cRe `�e�g�guhj-j!k  �n?oQo�o�o�op  p4pmp{p�p�p�p�p�  pnsvw�v�vovu�x|.z`(zz� �{v�z�~���� �������  ����������  n�~�~�~�~"~�};  }�|��a�つ�b�M�8 .�݀ƀ��܂P ��v�׆g���_�Q  �=��ň� �牯��  ���`�d�h�l�p�t�  �x�|��*�Ên��  �������󚤧  ���~���J�����\�O  �E�0�����v�*� ��  ���_�:�.�2�^�ŷ  ���������t�N�˻y  ��O��ȹ����e��  �����e�A�)�Ϳ��頿���"�  � �@� �= ���� �@�`��������� � �@�`ǀɠ����� � �@�`׀٠����� � �@�`������� � �@�`��������� !Aa�	���!Aa�����!!#A%a'�)�+�-�/�/3A5a7�9�;�=�?A!CAEaG���K�M�OQ!SAUa                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                MZ04   12t    ��R   !PKLITE Copr. 1990-91 PKWARE Inc. All Rights Reserved   �\ >      > �. /u                  ���k  ; s-  ����-% ��P�"3�W�D��˴	�2�!� Not enough memory$���S��9ڌ͋���������Ƌ���NN��+�+؎Ŏ�� ����u����� 3���� �7����A����B����H����M����S����g����h����i���r���Jt�s�3�3���Jt�����Jt��Ӏ�s(��Jt��Ӆ�t��Jt��Ӏ�r��Jt��Ӏ�w|.����3ۃ�t*��Jt�r#��Jt�����Jt�����Ju����Ӏ�s.��,���V��+���&��^�v���Ju����Ӏ�r���Ju����Ӏ�r���Ju����Ӂ�� ��뼀���Ju����Ӏ�r��Ju����Ӏ�wE.����t�[��Ȁ� <�s�N�P�� �����  ����Î��؋ރ���Î�X<�t)�������Ju����Ӏ�r��Ju�����.�����[���3�����Î����&�������Э�����S�P�Ŏ�3��؋ȋЋ�����      	
                    	
         :� 3�t���,��	 �  !"'(62K  `D9:;G<=>?@ACNOV �Z[hlWLEF  W�A �.� ��=��t x�w��� u��  �j��ȻUU���u� 	�H ��u��E�؋�u
y���u�.�J ��  c�u�� �.�q .�.��sQ�Fo��0�.�&G�C�9'��>�.�:96&�m@ ���Yu##t�.�&	��� ����`�)$������6�v�����	s�?HMY&�f>�2�	�AV t.M�@u1	 P�u�B7Hky�Z�g�.k愍�{:u�1�4��?����@�����R `Q UWVRQSP8 .�'<&) �.��Y
[]y�_6c>e �_a�gsxi`�3��R�Z�ۻl ��
6 ���O����\�)z���;{Q������E����}Q�����E䇎��&QO����.�����GU��ۗ�r���U:%=Hv���t�qP
@t]Aw!��#GL���a9@t�� �"s	� L�e) �> 
s� �RP�
]��QP'XZ��?P
  	���t}	r����t0p-'��� ��~���nI1�@Ig�I N� �PSQRVW 
�7 �K ��d� �� =�t��0 �(
�D/P Q����Y ����N ]_^ZY[X��S����lC�;�r�C�3P@=t�B���PP���CX�B���;P�a�aO	$�	8���,o	`t#�]�T��3�����%g�@��/r��Fp��v	pFaY��
�	� �X��:P� �����3�����d ��6����	�|����p"�.�
�N@��U��5P5P7FN9.�Z�3x��)1 ��.; Xt�.��&-� �3QVW3/�'+� ����>� �_^Y�H*$SR�#J.�>�t=��aZ[VQ�${�	Q�Q���5����>�cj'��m[Y���1��.+;���6�5��7 �]4���8�3�) X<w� �ϥS��\U�.U�f�U�� �"X�  ���9n u�~��t-��T��J�&�)D 	u���P=uG '�;�t麈a�<\���#; t&� =,	��" ��b3�(_��_{�X��a(�aD!cpc.����jB!��|TkA$��3b��uto���z0��&	��8�+u�l`�l�����2��=��0E.:&��u ���VDt��DXu��1I �»EH�ER�X��\LN<�����<�����c;�`��&��_�;^�U?@K= @@�HW���>�� jC	�	A	 ��> r�X�>l��V�E
`iXh@_.+�b8{ ϜPx� )t���-�  t%���/��tS.�@ &�[�ش.�E KÊJAA3A�+��A�5�?�G�YGm�r�c�K&��(��S�V�Z]j,�*��׻)Z)�)�PS.�^��M}�f�b�yh[��QWP��2K   �>��+ ��S�* +���W��u
� O���Xt_Y�x���?.+- g�VW� .�6A� �� +  � -��r3� s�`4 r)���r%�'-'+��'��'z ������_^�P8c06
 �  � ���I�< t<\t3<:u����   �t�1�zX�VWQPgRn @�?  �</u�\�
<ar<zw �$ߪ��XY_^�W< u�N����"�@WV-��;��#��=\u� O�YI��?�O&��B:���OG��VG�
���ti<6� <.u��C?t# t`�.t����&8��R ���@	/� G����R�}�8�"�8urR���f;Td5uX38�F�p��� 6��� �\����!t
WG_un��i.�8�"�9�2��@G
"���G� $%������^_	+3�#d� ��� .�� 8t�3	�	`>�u��r ��F�|:tH���\u�	 G��;<�7/� �P� PX� C<* u�> ��I���`���%t�-�y�����N�g�� 6�
�.l���W�*���Ò~v�?�8�=N��@ҹ	���@c �!x:\S��ENTRY
\CO�OL.FIL Pabcdefgh.MS ��" " �)!!CPS.*Vi'�6q-#A1B2Ct3D �"(6ܨ9<@�l, �=AC.�B���x�>H��uh��u�B_�ܸ
s�"ˀ��At~tpt>a�<tHlu��%L���F��`�>bg�6����u��8_�A�"v�R�r� �.r��r����	�rޑ	@0��-~2��nn9���	.tf�"sm� ��	R�s 	����s%�.�@�AWIs69�)� �$
s��[�����c�L�c���4�+QN|Z���&)bRbc�;"�<�|�j�<H)u/��ł�����R3�$��@2  �C2 �t߳�*�f��&n��v{�Ü���rk<v�z+
 �ڊ<�u�G
\O
���`2
 �v�og�Ds22#8��G�&�3 "_s�p_�>&E�X�6_��\� �� ����vm���e>!�8�� <=ux`
��� �<Cx��-�<luD���� /�]18�eu���$�<A��Zg(� s�	���A̤.A��tre�\t3	/t-NV�<v���6^r<�j�!d ���p&:uG������t3@�t uF��� p�>nVuqJ���oe�i�H��1	u@z���/sM4AUH �$5� �3�\#s�N ]��w�7t�ab��y!>4.aNh.���M�B�	 M1�� 5$c@2`�0�*hÜ��u(PS�Qh� q �>! �P����n*�3��V3�,!3D&!.� �l3" xHI$��nl 	�n�TX� pjr�<u$���*t�a+B�Q)r�2�����5>Z�1 Vr�HO$@_Xs�5�  -.�\��a�gL�tFl#��lr<Zw\t�'/�@�� ��g���xL1 ����HX�u<t��^8��^���p�zr%2�;	�%ht�}P��u&�E�\ⅈ�^�鱤��m�؉D��q	��՘Nс`?,z
WQ^�tv	 P:x.�c��X�!@�����۸:==�r�<�S���mf� �P�ظ	D��@3)8ҌXrF��z q@u?P,@���!�2�Xt)t2�A�una��У]e�G�_DH`�>�A�[,,t�0�@.I��@���,�7�CM4���n��ft�������;����ࣚ0� > ��6t�>����l��� $~<R���	:�v��PR�,A� ��7y ��=Ƥmr�ZXQ蚸������q�]C�����r3ҽ�� }��pM��7V>O�{@BQ��W�dV�4�_�Z�@� G3�F;X!�u�$���� t�Al)�l ��e{"�N=�K�YI$R??FM�NI�I���S�̄D�"
��h��o_�#�jd����Î[�U0t���(����!NN�q���Fa��� �O��� �(l�]^�,�ϰ �ԍe�� ��>f�.�����ri ]��߸ A�Ra�[bR���pdr�`�n�5��`0���;�r@���Z~��8��*��r
��V���ô9��Ð���?o?��C�& ����IH׭53(7� ��77���(r��x9s�B��;���`��.�-.�qμ�ht���r'v��'x�.�(q�w�8!x��"' :� W��Yu"��+ϋ�f�h�1�.��<z��g�ÕI�>�H���9��iP�i �d�\p��v�D  �uߨu��� r����rу|�� Pt;�ww7�9s&kVY �u	�L`�^Z�É�ݛU������ɔŀ�Lr��|�
��������y�
�Ô��VWQ��8�T*s�Vp��(+h
`\I�^u	ڕ��(�=� 3Y_^áYY �u� tW�|� _Bwqsr1�s�t��pDuA��y8��|��!�W/uG�9��]�s�ċ�[wJB f	�R� h.sȑ� ���PRW.�E�4 ��c6	�+	�	"< # �4�.:5t.;�u:UX�}�����_ZX��, �$TMPI0PMGTHMX �! @
W
0� H�_D��g���m!��� �R �����ÃV	
��&�ܐ.Gr
 ^(� v�Ddut�Lsr��m0Yo�s�2AP����u0	��F
Y�,������ӟoRx�*��0	�����p�m.�Xz{�Z{qwU��1+�{�G~N(�ub��9��I�� �|��Vՙ��jظ Cxns��QV�<� U�<Zt9u�A������1N��^Y�J�g�.ԡ>�8����>{�����;?��`w���ȣ6��>�'&u@�u^�6�!�^B0`N�,�y�D�i�?�:|<~YLp�t^.k�\Lt8.9 �t2R�n �C�Q��,I����RrF�7�Er2ΝŃBS@�� &#4�B��0C5����&�����sT�yO��C=��C�C���+P�r�	��`�r�� �	��|�e���i�S��ϰx]ZA	2.\d_
7	.�W�[�#uV#	=�w]��	w�+��|g`�H�Z3�t ����� �ʋ�i�6/-� $��2I$�0� �9����VQ�R `	N�^j�)��zw�$�F��Yz��ό�K'|��1�ͺ���;�������f.!�h�H�Kp� �-�����-���$�g �>6rw
�$� ����P����h�J�u�l�ˀ� �ue� `���ʊ���r�� p�.{�s�Ko:�+�{�Z�IQ�Dxuk��N���TR腆8M�蟸��dk�1��r^�#uV.�%$g �rI��<uC.��̌xh��I��(u������}�3���"IVI5s�G���:`�@uP���D@d@��p��� �»j�� R�
UoD[�����?���� ��jH�I�Dalu�$�z �� tPlX�0����LArZZwصU��A��,z s!��r9�y�G1')��Cr���S��p��K+�I�;s��  9��N� ���� �y �t��A�H���PT�����1d�`�
��~.cd!�e7�.����u{�u��6��.�>������1���H�����6�EQ6�6�1�E;�6�6_��6��Ն�+�v���X~��~/��6{�z�yǛ��viC7jt�k &��S�H2}�%�b��,�[$��>_ |���6$�N�6 ����2i�ӈ���*��鄢�@����ch3S����;�w�|�kbh;ց�̀�����j�}3!���1�c�]�!AfW�&YB<"���a�_b2M�[�u�Zc��rqBZc�Z�m�kr-��}���dV�6�A�z<���e�7R3	ٴ: Z��<t<u�O $19�t&@/�_��-M[��+�,�7�g��t$.*;@3v.+i�Us.)��p��N�,�,\�\U
訆� r��DE? I�8u�Zn08�S�1��6�<�H.�>������%	� �W��S����Lt��l�wL��
L/�L�%�L�n�������I���>W�7�Y#�9B"!W�����3���tP�A�� �[���������"��Eރ�]�	���r7��`���P����Xro�&��*���rc���,(�]�v�?����rD��?�Q�*��k���4)�j��I'�[� � ��[��fZ$rP�`��	�$f���-Jo2�̝���T�2��sWͣ�X�!*�-X�u�*� �F&9#�C � =�t�r��T�ش?�;�C�7(hu*���6� ����#�
�ia�PQ���N��� ڻ�{�W�w��lc��F&H��l� �H� �4�r}Dt^Fr/L+,C�Q�Dr  *� t�\r�os�����W!���a6���/�:�A1R9����f��&�*�+����/,0�% =u��@&�Rg�1�W|�VW����A�l��rck]m�S�gOe �ێÍ�&&m�&��5K�&��&�T�w�P�_��>P����u�dM �X�B	z[z���z��hjf
�f�]�n&�X�4#&v =w;�ƫ 9�W����h����V~�<Wz=��
�=�_��d��� M�������A�	 ��.��2���	�b��v Kqa��uKm 8s*��C�@�2��� P�9Ov����Ye��L�2����JH
	�`6 NJ"P�����Xy������t���� ��Xf,5�̈�5�5r��5rr22vqF2���z��̂}�?D�[��~����Yo��6�P
뀛P�}D*��/OZYX�^z�����PCTRACKR.DEL j�t[c�Ng� �'�m �˅���/`��u��At Bt:tL������	 ���O	�y�&J��._���R#�'}bŤtd�d@��� �s
.�H� �s�j @ u�P�'Ost���s�l�.Dn� �C
���
"訕�\�q��
3p�y�bHs	k�પ}��;T�\?TU���T**�h	sA��>������B.���
d B 6t �#� - .��!
�CG�
'G��OuK��I<�����ƏO�� ˗u, �$.����$���w�����_�%�K�emJ��&A�<� rF�u:�sY`���v/\3����so�1:~��^l~٬o:�s�=�*y� K&�>� �� P:~w� ��M� �G�1� �S��kf$��/jj�< ?� ���>GE��]u� ��iO 6��F/�p�E�W���(7� = ��w+e@w�AK�wj�2�w
 �9���rZ.�����B�u�L��Ft��	�s�=�v�2���
Ib f0s	,�	1�	$[�D�Vq������2��%�.�r�r#Y0��@XR�`CE���t	E��_��[Q�Ӎ���.�̀�.S�+����d�&Ρq��]�a �͕'L]q&!����r ]���ɁMu��T"� $��� �
GJ&��9x=n$5+o� �L`j]�م+�H�H��u��=� tt���kPR�M��@��i�.��M��ZXt���ƻ�0��]>7 ������T7�бʻI&��@�~����=��
�R�
�ѿr���r���a��.��Mm�.���{�@���������� '٧7�8ǧ��)��L�(< ����À�tQV��W�ώǋ�	����_^YR�إ��Z��z���!����.�. �)�j06�� wu��T r���{��I���!���5�:ݾG����rƠ�rr��e�Cuܗ�, m�xM�k��_�r��f~ _)�H�HH�>w8T�v�˧H�ޝ{�]�HS��ΞQ|5�d5�5��5�
��5��*$+V�x) I^�� ے�� �� �%�� y���	�P��-Q�	�݄�&
�$�&����O�\'� r=�|��
	8��yٍ�&��h6����� ���y:� �a>|re��>N\,ǿSt�%��K�k�� �[r<';c�8�l�u-�G��;�u#

�Ώ

�umc
u
�u��
>pZ�= �i=��sd�����YtTwJ�Q�F;�u�R�z@;wL1�84�&�EwJ��[ED!w �&�E����
륫�� z��6{;�s!&��t&9D�r`-v!�����t
۫�1+�6�0v^?t^��4�A��;O��Ȇ��$�CZ�T�_�7����� ۯ��O�� ��n�'�� ������P�\���uu��S�D��%�6r
����Ý����ILU��U���Uk�X�b2��k��C@���v�o	��)�r�s���˩<3���~E�A�8@u��(�� ��vXr!�	8�<�)9h���QVV� ��6�nx�΀n��}"֚"&"�^��t��PD+� A��F����X�(��[P.u���q*��+DP�w/$<@��6g ܋+�tW��b�_��+�tR�?��WV���&܈����1Y��a.9.t���*g0r#P���g��,�(c�,�*6��<��0_� !tf�]�(��7N�9���c }���n,$�t���%��^=��w'��}{ :�r�&� ��2�b�t�z^w����O�*)��:nuQ|���+Q2w=4�}8&w1L�
.
<������*�	�^_��d.��������	�!�Sa���t?r��I��u��A
����"��ȣ}YtQ���)Q�B) �	����!C�7�*���*�@���(��8(��$r ��#a(��G4� "�s �r�>  t���^G�JyO"'�@��<ar<zw, �_�� DATAMON  M�irror7�pOOLS= `CPoint Talk���t���7��SENTRM Y
\abcdefgh�h.MSCOrz.FIL �!�S *�/�k�MN��#A1B2C3Dl13
�����أK���#�� ��qY�ū� �mn��7?m&�'�1��>Jcx��\U��V�NZGap�@6��Ct�N��  ?�S�!5�!�������[u-;�u)$l�%`f$u�&f03
�/x@�u��� ��=��	ڀ�z�J&���#%}�T���	�� �#�y����.����uh@a��>��9zIj���y��|6���� &�Y��V�7oX�W�<�Z�[��.�ڀ�>��Ju(�q�2g�q��wt�6�fRP�Ģ�XZ������o��h$ �a�Z	�S���L!E6�1�\
`4�R[��8�a$�V�=�Z�3
�A�)&�E �r&&�6N;pр�r(���X@r.�p��Xx0&�&�I��K�r#�
x1�H���-�O��/l߾9��!>�t8	�Z,�z� 3�3�ɸ�g��UUu
;�u�{�Fy��ͫ���s���ii�ؾz�(��*�>4�����7>0�zt��.�	H`��)������Ѣ�6�#L� ��@�!�tø�y=�2~��	.$W�%e�VX�&z�Z\/2��4�  �U��0��	���]	�`&�	l;%��Q	3
}"M	�@&A&EtNL'&�.#��&z� ��E!���b��9�!����8I��S	y,	�J"��?u�#�R	@u�e`�B��z��
�&� &����8�����
�� �J��;�t�-B .���O�N#SU�!!8^��&+� ��VW��b�O���6? `O�t3���$Y@�[��V� ޻ �VD�DX�1I���/�� ����EHu��ERu��1 "u	�& ���0� s9���=u���^�30�r��r��iF��0��eG$�Ց '��	/�ݰ� ���Hذ��.�&2rj.�ە(,��@�y-u�����M��������D?���7$<��W�4�<u	��u��� ��]�O��k�����9� @^�_�y�W}�7VN��3J���.20/�/���/���/���*���A{ �(��� �� ���k�
��C��}�O'�B� � ���q��N�.� K�Bv����A�.���D��/�Q,@�crG�/R`�yR�W�5�1+��/Џ�#��E[�O� r �r� ���d�w��+'��UE$+�3�3�_��L���o(��J�l6(6��>�83�sX;�'7s�R�9fxs1�3w��n���v��Ó3��t��rA��# �����������#��'��}��x��OG����� |�� �	�<��O/�0\� W(�6e �p< t�\7���SG _���>� s��_��ű_�un �"4�m� ��O
8��Pvy �_� Y�r��*��Q´2���f�N6�_2�6B�DUHR�*?�:�#^'� #��+ ]��ʠO��� O��������F^~���$Yo0��Wt| �+|8��D-��@!� S4���B�O؍6ב� �� ġ�� �$QW 0���_Yt j���WQ�� ��Y_�Ç7�q88r78�8?;0��0��)QVT>cD�|��A	^Y��~��5�~�(����O�� ���� ��	�� ���zt��� H�� ��;�!���  �ۊ�� ��ۇ�����t��v���/O,�,5��f�U5Y��5rU22���2B�rF�^/�;.l�G�o�w���#'�? r"M$��W�DE���(h	��Shha�<�y+�qWQ�����Ŏ�����w�'P�����NI)3�3�&�9{G���ǌ[�����9��+���\��%�	. "K��2���.t		�� �� ��!W Ԣ�a"Ba@� ����� ���)��� a�%� ���+x.�I9�$�'ʃn�A`���sC��.9 �!s���ڶ$�r���	���;`rC� ������J�"��ψ&��E��3�����&;�5u]��"���|V���ٌ��Ě�+B����CY�C
��C_���'�R���BoW�� �3��1�s���O���@�! ��?� u��;?���p$� �tD/�<Zt x<Mu6B&W�=�=��,`jtW'�`.&�u�pVSCt�����dP�[������r����Xs�`�*EI�Ɗ+��A%t� ��;�u�(����`W.�>n� _n�Rl�.�SN��&q�O��t�.Z��K  �; r/܉��6^`�>bGRd�3� ��!;ϼ�����6������u��&�G�"��B>&�=&�f��/Wש�_tK�G�"w�6E�_�D��1��	Aw�wv��Initia@6lizing   � control file  driv	x.
:�$ ��T�C��� ��	*Q��x�525�0f�	�+�.�p�!,.����g�!�$Q�r[�r	]�l�s��@�<d �A�g4�:g\�
6I�_�f�S�� '�2��z�p�E+�f-�t� >�%�������=1��.�z��� 3҄��B�ۄ� �tID~�J�DI;�	t8�:��+3��$���th�^�//}&��B�V8�8�% r�$r��,�p��2�/ ��3���r@�ۅ�8M<�{l	�d"��£���������'�4���۝��CrU.��CxIr�F��i`O�&8�8���nk"[]�&�#�uv�#X()L��53@��� X)�	#+g���B�4$�)Y8�� �C��Ξ��'&�����6e�s�\Y 1�?U�0�3ŷ�S�+ u��
�mAr����x?���B $	��{�.��h�ڸ Cׂ���� O���:�bD����r7�����r'�1�y�__�Yx�D\r�� ��
�G��+� ���G�p��=v�l��@ �M)�,��sWV�8��X�'�6�'.�6�?��w�-���'#�?	�'�qb�c��yc�L40o�'�M6����3 �t2�l\H� 
�'S�
iRR̨ 
�'A7/��7�7�M1�u�^Mc�L�L^��_Q��čB<ޫ�-�-R\� ��-�1��� �k3������0���� ���u3Í��+w<Ǽ�}���'K���P+P52���SS�H�S�,��`p �[��3�)u`� ��'+��kyCk]npn�2��<n%�2k�1�2rW�!���8��t�΀t��2��*��7H]�+ u� ���.,\F �O�wr$����: u"��:�\i:zPr`P i\*X��Q<Yt�{<Nu���0�s=�M5s_��&X@$�6*��IP�4@��OJ�	��4`@�<J�O�s��64�;2;�);�����#B	�7s�LtS��?[����`	�������ǖ� -��1-;��É$3�����S�`�z�Bz!�; ��u;�u.���̴YPK�>���/�/-�\=
[� LfiguratÝi
]�[ �naults][mS�.^ [seUUwy@C��  arch=days=p{eagslo�AwV$t d. n6=ack%=� Fuf e �l TRUEFA��LSE54[5�<�e �Z!�1 	�*.* -TMP��VM?WOAH�SWSPL�(RMGIGDTHMDOVGb'MS��ESd=P 0H=\UNDELETEj�uNI v����*NoU�+ �����]M�>���t܎��C�>9kܐ4	u�i��� ø� N� �!W�_� sh\�	 ��YI+� D+�+���p��
�&9E�\!� QWF��6�	  �t_Y��XY��;2` �&8t
%tG����Z���T��B�*
��"|:\uC�u�K
�/�!�.��
Bq
���2�G`�
f�� Y�I
�S}
��A8��A.��	�'�#t�_�n���;J�j���%�G���������0
 a�\��'a(G��
�l�w
Q�YY)"�@�ZD`���3����
 �dZ�D��Z�	��ZX��HZ�� \��� s1z������yxQDc�ػ�YK 7GMG�1��U.�� �	��:������<\t@���&�}�\uO4���: �	����9k��E�y�PvZ@��r�@��w�[�&0UO=�Q\ڣ$$  �
!� r<[u�������d��P�*j$��?"<C'�rB=u=�'�pD@u����  �<	t�<
t�.:+ �t�<Ar
<Zw .��-�&-�7����z	���f�<� �/F�:u2��~<]u�DkżÁ�Z?jv�|��.�;rp���F��?���F�R��i2�t-@	�g�]����� �LLz{�1&R")�I�Y� Qu�NP�X�� 'u)���'5� v�Lu�1U��11�U�1d1d��1�1'���2� ���t�(��c(��#���29��cP�z*��ɭ����X������y��u	0�< u̴���X�Xkr?X�6ӄ�Vu3�!4W�M�>�2�{ĐF<;� u;W7;;���a�zP�DR�[=�2�� ��a��.Ǉ)�w&,&7�S	���ur��.h%��C>$�T"'��� �r/<t+<0r-<9w)ғ�u< B% .�
���
�9�Z
��<���
��W�����	�!�		 Å��;��!S�F�wy,�tc��u� l��t�F.��v,��\��� <	E��/�q�����7�z�H����W��}	��5�	3��	&�&݋TQ�譏0�2��2�����H)� #�U#��o��R�1�1^ *Lm>rsZ:��[rg�n rb��J!V�g��QjafE��@?f�
�4h�M�� 0� <w�t�=�	�!sSA*
)Pd��� *�>a��>�
C- 
 �'�A�Q&�=�
�t1�IOr2,�m�&�P�� �33-}8���5Y⁼� �|�(` =c w	BI=	�f�@l�&H7F����v� �ڀ?^;�v�r$BP����k?���8����7�o�d���WVU ��3ҋ��O�'�������p��v�8�������0�O�<�'���'� ��]^_qT� 

�
 - A *LS proc� � facili ty)Copyright (�AC) 1987-93 C��al Poi  	 Software, Inc�R. 7Al7�seserved��TRtod�p�revouslyۄd wvh ��
��mma��n:�[[��7:][pa�p)]Jname�V/DT | S�OS]�"6/LISALL@PURGE[DRIVE]RATU:��LOAD<S/
D �V/;��T-���]y7�'sL�is��av�6aab��to bre��r�8 �^�R#N  ;out�mpa�t�for �#�rm��KC�Kl꥚as���by MS-;��D�^0DO�Q<DcT֕.:eDSDS]��a�^��Qaoad:Un�֟o m,Aemo4o��tJڝ�DleLfZL�16E�*�]6PPurg�ll.cł����i��tIv~Disp�-lay=�����d�OVeff!;�eachʞ�P�@�En_=Ks�Oz�ofTRAD[�}&]D��joCF81�, � �FORM� :W;�cSpXifiv2�(x:�m -ja n�work��N�: You c�yyڊ�cuse����
*7Qs�CKۍn$$דat0pRySUB��aw%%�xZ��������T(e�'���.|*.
D�]: F���=cD�s�{Invv��p�@��ڠs%5?�L"mhA����K.$Ni�7ne'Os mutu6exclusZ3#x�c�8/����0���0�-t_�#��f�?ou(:U�w�s!�. B
a���r���1�AI�O1B'#%��,y�+�1v9s`
�;u�����ԯaD�.s'0�g�@�����<Of�os�L�#	8_haFHncPswKm^,�v57s띇e8Z>6�̗9�*�YH��[HPE)"*g"	d���/�o(�Re[i�D��k:9:{g�8�ku<>�-9tC�B�4IlunB���`��/G��Us`M2�0�H��={'(h��$���'I��C�.ې�
�Q����Insuf_	�Vg�ua�]0��|$NoB�e����Ty԰����$2Fc��>]��6R(��!�=H |$O�����+U�t|Μ9 D�y���w�tojk�1��5c��VU�m`? (Y/N) �9�n}q�T綜P���nzk	�eo�/�A��Tp�?7D�z8)100%O��H1gIuStU�H�7Y�4���"��S� � _e�C�˄ p� �SENzTRY�1I�<x4H�Mam6ype�ihdc��H*S��"�fAI��atLB%B���=�9��;q�n�&-�^an,ړpV T��;a�� �r�:�*qFI�5(a�1%A����z�z�)G�DHIg�Y�e���succ��fu*�,���Ood�Y0&�<9. �Aabo��r{r Ri0�3  $���@������   %%(%^%r%� �%*�% ��%� �+&G&	a&  �&�& �&@�&��&��  &�'� '�2'�H'�U' ��a'�x'*�'F�� P�ϫ�Bhy.8eft,�cr�FIpLES= �u� CONG.,�SYS6Va�n�*% ț�O%�'co)E�rK x2�+~k�wn)�$U
 e/gg B��$ �4dis�$kdؕY!��%}�.Ԭ%8q}�teHn�<w"t^K�a��Qe&@�0RequeK�3sZDMA ��Vruf5X=4� Ab�W%�ZǕ�64Kfw�;a� MȴTia 5"T�CRC�O9�'�C��Bl��u9 Se��ekte�WNp��A����P))�dr��cam�[�\�Pr��І�$QaxWH�<�/*W�UnI��pH;1�%��t.t':�� �C��
 %Ҿd:W�1  ����Jld��-�ylN+A٩�hG�Di�]Zt+�BPCSHELLN@0DESKTOP'�0COMMUTEC0BAC`ALK'�1nee	�op4?s	c���/(	u}/�2WW"ows	�a [ta���sWch�)WBpm�2Gg�MON0�5�._K��Y3��z�la�Ast7]7g�,�O,s#mb�ryROD/��&��_Pg�2g��
�A TSR�nks;� ,x��|0$X�%-�E��~P!Mb�Z�$#�.�f$}Z$NONE6�d�dZt�* \A,�c�	� .,��o� @ h�|+u� ��$� N�@*~'E-QX :\#%&-012345  6789ABCDEFGHIJKL �MNOPQRSTUVWXYZW�$.���!.#$\'()��-@�|!@kt�^_` {.}~N��x�PCTRS��R.:л C�	��*.* -TMP��VM?WOAH�SWSPL�(RMGIGDTHMDOV' %�3��ǻ �� ��/���t�=/PW���  \+� 8�!3�S.�&G+��6$G� ���������r=/�ϔ .��+��g`��"��.�> �;��9%+�3�!�8�͋�g�.� �!.�X t��	@n �8��?�ȑp �:,@tc0	�t  �� %L2u��� �7��{��!�i}6�t
.�1��%Դ}B���(��S!.�!,.�s" �EH"�$�5'r�(� �<Nt�� 9����.�E+*V�f-�=-Hr���f-!n���!w%��-���)x�e� ��.�q��sռ �;�t,�R�=.��L���Lq_��-�
��t�:5@�U�T 57�)��=���1�&5�&P�����tS .��+&�[,V&X%��)��)��)/lR//+��;� �>.,� �F ��O.�>P/}�\t70&�\*E.�EH �N:�/�G o�{.B�Z�s���?+��� ��rU.x�.�+j-�݀�>�u/�r*  ��t#� u�Nr<�.�(� �;r8-xd6�����;.�+r�`F���6�}&��Zd]"�� r9r]]���r
��*Ā Pă�y�X��<�(u�����;p��p3&��Rp.p'c�p �pmMB� �ц@ �u�`q]qVWQ3���W��t����Y_^��F��'X�	
A�|�' t"d"�L��� 	�f#$r=��P��x,  ��t	2���# �	6"�����#r�P'��X�V%�F<Nu�?�Ǽ��lw=s-x���b1�>���>�>�=��0E�ͼo��ơ �v��+3  �����������t@ .�C-�<r
92$�d?��j
S
Z��аWV��C���-� ��>�-�^_�vb�3n�~̌�%��O/#�܂��m�< t�a�d�'����S� ��.��z,[p?��VRȹ�cFcO�= u8O��g?G�V�װ.��  ;��G�:�� $�Z^�p S<�r�[+v �$�S��`�[<@.�[������yx6�&Ղ��p&�\G�b�j� \ C q�!s= t	S���[����A�YC`s5.�RO]� f����� ��s�+�tP)cE&Tw�� 0��+�N!X�җ@��.t@�K- � �#s�� ���3��.�. .���T!DP0�-�}���P���Q�#���ީ� U��C
�����f@�s�93Tku\��p� rT�ŗ7!;�C�PR�� �ZX	��)’��� r�@�>�",�0"r�
����PSQA�+�+�� ��+�8;���P�='�ͣ�����+�� ~s
X�.�3��/�+X�� ���ZY[�X�ZW.;E-sTcp c��� �@!C����0g@�>t
�u	 @�H���|��_i П�'� ��x�� .��'.�33�"�'��8	�'?+9N?$3}��̍�'u��j�xu�'� �Q� �t�~�tTvH�t&
�'S��uR�R� 
�'A��\��s�**Jv^6��1 �"	
���j-F@�}T����8�9w��6�.��P���&��� !��-.�����-�5�J�-hWjw� _�%�%����!nr]񐂶-0u:�t2��P=r(� 1H�� r4@���.�h-t&a���G�K@p��)u=�8hH�����t�O� m� t�'R��-���Zux���R�QN�����5I�D7����tX � �}�x�����rL��X�@�xn� ��C������\u'�!��G�)�B�ܐB�B��%�u�7�X s9�st�\$�\QB#�23#w�? �
�f���� ��@s��"�E�I-�ȈG-��h>D.#@:-�.�?��;/�C�&T-�(��WVhr-�	[�-�A^ _&�DP.� &��MD.��-�4��D���n	r��n�[=9�	v�b���|jz��0/�G���#������ uC.��tV���L�=#""H��ʠ� �g&0�E)A��Vs?[�|�~^u�sㆹ�}ζ-�O�W���I��6��2J$P�7���k�`�R`ԡ��E�U��s�>�3a����
�_ K��
�`�l��À<  �7� F���QR�I9�
�)���8�!w���� �
[���?ZY�E�b-K�V2���� s�H���
]������7#��>�9E�#��->�X&� (�x� rs��?tum�fu%4]t�{d���r_�.t<�,���O����c�A�2�-���0��u(�0���A$��  �� ���ʱ�
������0�$r����4����,��X+3��/g� J ��)<t+<tP<	�<t
��� �s.����Y G.�C�5����9����� I�/u���Kt�M�u98� �v�O��;�P�.�;�P���P�o�P�X�%3�
8f�PQS΀�-�<I��	[���˙��$�Z[YX,�S��vDCA �6&;Y��  E�.�."`��s�Xp^�+��!�8pwP�s�+��B���+����?�0��=S�C�-QW  F�_Yt�� �p��E�����R�L��EU�N-�bN?�	aھn��Dj�$UDr�d8���+���&�R&C `-;Twr;Dw��1��d�-� &��+k1O��k��wt��R��i�$$
���!�����.	��: %�_�P{m
�X	I�ăOS4&C-��,��#[�H!���[�K�20��:���(�.rL�"�)` �!���Zr訄���h�,�ڝu�� ҫ�s-�a���}���m� ��ī���>$�� ��/~)�B�L�-D��o�$y���D�-�b�.�I��������7�7�7�{�B�� �?,���Φ�C1Y2P��k�6*U�6�1����/���(,uF���PQBFP*.�h�iy�L�2���{˵4�{�c6��^K)(7���Æ���"s��Bu�:�r=A:�:�r� rt��$����H�Æ�$bK��ѷ�WV-�_�� s� 	e@��E��E�?<�HQbt}#�_��_.%�_륟H^�%М��h���u�FS9N���%@��t1��t��`4+�ʊ/�ӭ6-��D�2-@oWRV�h�\�kx���,�'�L�S[{�)�t;^Z_[b����l�p�$�	������d ��� �@�� ��oʋ�.��Bˉ�˻*��! t	$E5�Q@u�!�@�#]Eud�㩀�]� jTjI6.PAi iyOl���D�\����m��F ��+���9'P�>�|>�-ON���\�$,�ny-�7��:t& !+���X;�u �OU���IFG�u	�a�lR$�{������RӁ!5#,�=?��*u��w������S���L�BT��*U�P�r�G�*t(IG�	Q!&Rު&R�R�$V �B��\g� �x��?�^u��Q�@WUZ ��S�Ǎ�$.׳���B.r���#ܞ��d��U귃�N+X�[YZ^_].�&�%.��$�@�VW��u^\�0�$�t��u�$���  8't.�?  *t�����Ĵ �.�p��%"�B�_i $�����  r�=<At<Rt;�맮����&P|t#���E��_^��
��l,l� a���	���X������H"�",�´2�D<0�� G��+�G���.��+�2��(���3���r����%��7[G	�,**���$����H=�v��:AC!G�q��+�!y����&f�s2�Tn�'����	�Bf=LI��.jR%�d����Zo�.�^��k�i�7�i�����f���#E�&zj��BBP�e��)�۳+X��%�4�R;��	r��]��=A��Γw�[�=�}�I�+	L���d;�;挻=�K�.vP�Hҋ6�+���+�M @�����r2H
12��<r_~Ocpa���ǎ����(_�+��N���!�+���HM��4�H�r���y��r?�����RP��2�XZfq&I�'�f{� s(�� �M�� �w�n���  �</td<Ar#<Zw����:u���.�px.�3 .Ah.,���!z:A�l��/,:�%m  X63�.��0,GFI��DwtkPr��?�P=4\�GT
1,^���caǟ�'Fg �K+���r ��=/uGI��6�o���=D *Tu �e*�n��u3 g0@�빈�%Su'%�%����u.�� %$����冋�,Ou(0L�v<6��z3�q��uۛ3X 43�h�`�=LIu)-IÉSTt��H�F/W���.b.�2�~.AL#?#G1^�T*-*-��[���8���C�t%  ��=PO4UL� Y�̀RGt���<EWN�5$�H��9�hh�鶏��b! ���x���Ar��_Zw�.�&&}�'(��R=RE��a��A��-�UN��u?�"LOD�F��AD�8��e�4-����u9�����t�����I�<Uu-��)�z)) w����(����������ou1z�l"l��lz�C��\�C�C@ѩ�lx(lе  �;	p�2 u���. �H ��X�M��-t��%Yh�(��`����(1�U�q��2���A��_���"r�K�ǋ96�H�>',
 yQ +�
��E"��r �"p���.��.���C�����<S��Z��P� �2=TAXtX�ܓ�!��{��`�J��ţ�ś�ԇ�� ����(;�^��zz��Z��-�gd�iON�7�\��#T�T�Cwʁ��"N���p��V)p�b��rp@�	D0�� u&�u�\8嫖}�:���t,�6�� �*sG'w�  �;�)�����0��
���
& B@t���_��c�=t�0n|",&�Iu��k^� ����<0 Lr$<9w P2�$�R �q�
��s�	Z*&��XY�����+u �mV��� �ށz����� ��fwMtg,t	t0�GI��=��<f[�À�"3o",�#l',�/aF/�VWQbr*���s�+ jd�+\�Ѐ�@�%i�+�h��  @�&��j&�G���;q�mF� ��\�pρ�/,��G�W7\uG�LR� _�w�:[�� A?�$S$0��rl�粑Y_`���{��\�-\.��#,�ׂ�e��G�$�"$	 + ���QI��&��f{�H��1��*,�X uN�g.�U*o ���, ����~.�%L[�[
���� Y���S 7 ��PR�д[f6Xs <�2��"�/�u�h�tHt�^u�S�s�ߢ �����O�.�'_����΃�vp}���y @E��0�O��@Jt
�����aO����o���:����� ����4� � ���g��+�AEX��  k�+u���	 ����;����z��^��Ƌ�J*.�.9%�. 41-�k1.���.�g%��3��h�2�y ��B&�X%?�!�<4���^\�ƜxG ��e�a= r-@p��gc�c*  SQM����丏������N���L+\WVU�R2$�]^_�.����	����H�=b.�R+p�����e}�3a����r�����0j�Z��+l.��P� p)r2��*r��}�x������ ܹl )���t@<.�55���*]9$U��I�[�WQL�	�	#	�FB�*c4�.)�����8� ���w..�����y�}�l�9 ���+�'���>p� �'�؃>��#e	ru���/r�C
<���;<�>1��La�7�c�8�b�E���^��w�U	�����l��J����RBN=B��r��NQ��.��r�:zs�V��*�|�I�+tZn�98��+tN�,�I�+r%PU�e�ϓ9��;�+"FC�Â�Ҕ����� �� tf��u;;��?;�N3�� ������= Sa=�tw(�Գ� ;Q��7 �b�tbw������*)߯�cV�{�J)P8wC�
6��,w7
.
:�]¿~��_&���^�a�+��n��8�N0���PQR�p 6�+��)�+tG0r��Iu��?nA
s�8�*x��x�"��Q#`uj��-H�hH� Z��]U���T����C��9�]D���+l9ls;��w�4X~�3Mu�&2/�]�N��@�2��t�|
���\�!���� ]Bp���V&q ϟ E��.��b+�l���n X�(��"��n��U1ͨC�(�9rtT��ϡv�z�:��{��%r�>ɲa]]V ==t?�D�� ���r���S�a��]�toBro��+6��vXv^�&r#k��MItsݦ�l.�u�����`}� }���u<ar<zw	$���n+ôI���p�.�� �&�7
��� �X>���� �9�\��>��>g�tC 9��� ����A� ��Y�
Y�~��uY�p
X �*����S��P�>��!X�Xи 1@j�� re$8d�6#�
=h=�׌��)�����	�'�x	�	/(3è�%_u3�u���u`2a sfD�	F2�	�(�33=	�	�4	3�	�	+	��U ����@Ȕ�u' &�2����&Ǉ �&�r
	|u�"0a��b��l���/����K
�q ��tG���rB��& ��� `t?��F�q @t�ɉ
 �x
]y ��sw�󥰁wm�*�z�7��r�H�d��)*�t+rov�+�J"&C�p-?��P:-��=�������B!����/
��q���uC�	<e��F�<�I�� ف�����  K O      B    Y��y��������!9l��������u���+S}��(7����`+p+Y�Y�Y�Y�Y�Y�Y�Y�Z�Z[ > u /t not loaded
  R6001
- null pointer assignment
 ���                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         ���� �,7MTMIDE01         MITSUMI ATAPI DRIVERCopyright (C) MITSUMI ELECTRIC CO.,LTD. 1994,1995,1996.All rights reserved.`+&&S&&&M&&&&qPP&&:&:���&&+&&&&&&&                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    �       �                         0	                                              �                  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            ����   ��      �      �.� .� ˜fPSQRVWU�Ȏ��\  �{�*������&����м����� < t��� &�G
�u�&z &�G@: rH�/���؊G�b�W��T��� �'�s�e$�
��y��m2��� &�G�z <v<�r@<�<�� ,������$�\��8�\��3�\��+�\�� �\���\���\���\����f�\ �� � �\&�G�  �v���&����]_^ZY[fX��&�&�G��v�����������`&&�d�p�3������������������G �G��p�&��`�����`�G��Q�= )t��`�= (����3��������������^ �[��� �a�^s= )t�w���^ �_ �2��� �8�^�_s
= )t�= (t�������V�>T� &�=������������U�G�G�G�� ������E�E��W�6T� �_��E�%�e�e�e�>a t �E�e�t
�u
�e�e�%��E�%�e�s= )�{�= (����{�l����������� �� �I����G �G�Gs�w���\�������������&�&�G��v������V�>T������u��&&�&(���RU�&�  &�M��&�<�|��ࢅ���>T�������&�E&�U�j�����Z�G�G�s= )t�= (���{u����W���>T������L� �&�G&� G&�G&� ���  �B���C�G �G��G �G �G	 �4r�>`�t�>`tV���Q����Z�G*�G�s	�{u����������<qu���<pu�� ���u
���` ��`�ʹ�>T��&�3�&�E� �n��>�t�>�u�6�� �i��I�&�E0	&�=�+�t&�E �0������&�&�U��&���O���C�G �G��G �G �G	 �As!= )t=u	�{u���= :���= (t��>��t�>f�t�>T&����L�f ���2�>��u�7�>T��&���&�E�����&�E&�U�~���&������ �&�:&��"��~�s= (�;��{u��2��>T���W��G
��&�E&�U�G$��&�E�"�����{�>T����������
��
Ī��V���������2��^��������������b�
���B�G@�G�G�
s= (���=����{u�����
s
= (�i��v����|u�\ �D�u�>T�
 2�����z��>T�D�����	� �,0����,0
Ī��,0���� ��J����t= )t�= (���= :���\��*��>T&�  �>�u&� ������������������>�uS��^[�>�u���&�G<�����&�G&�W&����u��-� �� �r������>� t%�� u��|;�w;�w������&����&�G��z��&�G��&�G��&�G��&�G����  �>t�&�'�{�����>uG�>�t@��;u	��;t.�6�����s= :���= )t= (��������6*�* ��*��������W���G�� �>� t�>� t����>� u	�>�t�2���>�t�����ĉG��G���>� t�G	���G	���(�����ĉG�>�u�0	�3ҡ�� �>� t�0	��s�������hs = :���= )�.�= (����{������>!u�>gu
�>%t��>������ǃ������Ўǃ����q��B����C���  ���v�� �>� t��)�n	��>�ul�>i�udW3��ǻ�2���/���u�J�>�
� �_W�OO����>� t��0���]� �s�j�u�_���� �_� �i3ۀ>� u-�� t'�>�u���u�ٹ �K���ًف� ����ٹ ��> u�m��m���u�Iu���t������> u �>b t	���������w��u�u�>�t'��t[�> ������~= :�K��{����@������>�����;�t#���� ���^�3������ ����>�u�������������� �3�����������������)����������W���G�>� t�G	���G	�s= :���= )t�= (�w��{u��~�3����������������������>�uS�
�^[�>�u�N�&��M�&�G&�Wu�����X������ �� ����PR�\����ZX;����r;�����u=� rR-� �� �����4���+������W���G�)s= :���= )t�= (����{u����)�?�K���������G�G���ĉG�G�G �G	��s!= dt= :�Z�= )t�= (�>��{u��E�3�������������������P���
S���^[�>���&���&�G&�Wu�����'������ �� ����PR�+����ZX;����r;����&�G&�W������s������
���������G���G���ĉG���G���ĉG��s= (�_��{u��f����� �\ ������e���	�>� u3��������������D��� ���n��K�u� ����������ࣛ�����	�>� ������� �\ �&���K�G�(�����S�i�i �k�k�m�m�o�o�q�q�s�s�u�u�w�w�y�y�>�uG�>i�u?3��ǻ�2���/���u�+�@��>�
� �s�	�u�\��?�� [ÊG.���G���G���G���G���G���G���G���G���G���G���G���G ���G"���G,���G-���^�_�G�`�G�d�G�f�G�g�G	� �G
��G��G$��G&��S�����G.���G���G���G���G���G���G���G���G���G���G���G���G ���G"���G,���G-�`�G�f�G�g�G��G��G$��G&�>t�s�e�>�u-�>i�u%3��ǻ�2���/���u��>�
� �� [��3��*���À>b t*��"b��!$��!��� �>i�u�@ �ػ� � �q�� �q���؊��B���w���>du�6|�|�%��|s�c�cr^�� �o�$<t	�qKu���G�i��� ��o��>b t� �-�@�Us�>�Ct��Ku����'r�u�t	�������ÿ��  �ra�q��B���0	P�tL���i��> u�m�m���u�Iu���>b t�� r�� r�u�t���	�u�����þ�3�;�sP�q��B���0	?�t;���i��o��>b t�j r#��b r�u�t�+���u�;�u���������u�@쨀t�=���w��u�@쨀t�%���Ëu�f�u������S��|�>i�u�@ �ػ� �? u���u��������u�������� �>i�u�@ �ػ� � �[���u� ��>)t�@�u<
�t8���w���^ �_ ����� ���^�_s
= )t�= (t��) û� �o�$<t�LKu���u�$�<t�9Ku����0�����G�2�s	�������&������&���������� �� t��������C���O�~�g�G��G��G	���s= )t�= (�M�=�V��{u��M����F�ð ���~�������G���G���W��G
���Q�����@� �~�� �u����G���G���� 8�t���G���W��G
�ࣽ���� ��  �>�uu��������������W���G�G�G	���s= (�u�=�~��{u��u����n�>�u�>���� �	�>���� ���� ������Z�G�G��s= (��=�"��{u����Y����� �>�t�>�u>���6�� �.�rr�F����G�G �G�G �G �G�G �4��L�>tE�����r:�����U�G�G�G�� ������E�E �(�E���r�+��������B���G�G@�G�G���s= )t�= (�8�=�A��{u��8��x��1���^ �{�����B�G�G��s=u6�{u��.�C�r)3��>�u�\ ��� �>�t���������� �= )t= :t= (uC�>tPS�����[XP3��������������>_u�Т��f�����XÀ>^tÀ�u= t!�\���=u� P����À��� �>{w� =	u
P� ����X�>tq=0tl= Wtg�>' t�'�Z�>� tR�>�t5�>at5�>� t:PS�� �+��[Xs)��  t#�� $u����a��� PS��[X�= uX��= Wu	�\����>u��u���= !u�r�= du� &��u�&������=Su�~��\����\��|�SW�������%��s= )t�= (�%�=�.��{u��%��e���>��u���_[��o����Z�G*�G�m�s	�{u�����1�����<qu����<K����<����d�������S�؊±<��ǀ� �K ��2�Ã� [ù���K����S�Z�X.������ ���u�u��u�[À>!�� �>g�� �>�u03��ǻ�2���/���u�|�>�
�>������
 �rb��^�&�&�W��� �>� t�0	��r?&��r8&�G&�G &�G��"� и �BB��BB��BB��m����%���$�% À>!u%�>gu�>$u�"� �BB��JJ��Ü�>!�� �>g�� �>$�� �$ �m� �"� �3��BB�$<tH�u쨀�� �g �w���O��^ �_ ����� ���^�_sU= )t�= (t��I�u�u@�>�u93��ǻ�2���/���t'�>�
�>���������� ����� ��Ê^Q�^ ����������G��Y�^�.��.��.��.����.�>� �� P� �䠨tX.�h�� �.��� �tX.�htp�.���p�tX.�ht[�.���[�tX.�htF�.���F�@tX.�h@t1�.���1X.�h�t �.��� PR.���.�u� �� ZX�P� �� X�Ϝ.�>t��u=u.�� �=u.���.�.���	���?@��
�g�b	��63�S�늇�6�b[���6����������6��
��� � �
�s7�
����6�7�u
��6��6���
��?�m
�G.����7< t��7�P
��?�T
�G�д��t�������j
��?�:
��7�*
�G�<
�>�6�t��7� t��7�
��?�
��/��| ��>a t��7��	�z �.��� �>�6 t/�h��(�g7��	� �� &�G  &�O&�G �\���� s� �`+&�G&�O��>!�t~����rv�� vp�tl�  f�� ����sfAf��� u��N���	�  �rC�� t=����"�!�`+��S�� ���[���sB��� �`+��&�G&�O����! ð/�5�!���2+�/�%�!�QS��6 �{��6 �s�$���6
��y��m2���| �� rm�| ��Irb��6��6��6�/���ؠd�G�`�G�a�G��6��b�G�i�G�G	 =�t�G	=pt�g �g�G��G
����G�>�6t�{��6�}��U��s�$� �>�6 u6[S��3������6��4��� :Et
��������]��T&�&�W[Y�[YÀ>b t*��"b��!$��!��� �>i�u�@ �ػ� � ��6��7�� �w��6�>b t	����� ������ ��� �u��� ��� �i��> u�m��m���u�Iu���u� �t�����J�>�6�u�>�6 uZ�b���6�O��<�u*��$`< u�d��d �5�t�g�'�g � �>�6�u��6��7��{t	�X �%��(��àb h��6h����>�6t3�*7��� �u$��<Gt<Kt<Jt<Pt<Bu��<4r��6�Ëw��� �� ���u�@쨀t�����ù ����������$��rC�o�r>�z��>�6 t�*7��� �u%�>�6�t �i����`�G�i�s= (t�= )t������ &�w&�F< t<
tH<tD<^t@����G<$t4</u�GG$�<Lu��0 r��C7���O7���[7���6���?�úC7��O7�Ê$ߊ�G�$߀}$u/3�=SUt*��=RFt"��=PSt��=TIt��=RGt
��=PJt�É�6�� &�w&�F< t<
�� <�� <^�� �����G<$�� </t� �GG$�<Du���<Uu�rz��<Au�ro��<Pu�rd�<Nu�q rY�<Tu�rN�<Iu�arC�<Vu�	r8�<Su�r-�<Bu��r"�z�<Ru� r�n�<Fu�� r
�b�<Lu�[��[7���6���?��F��OOW�
 �<$t$߈G��=$t_�5_VW�17�
 �u
�_^�_�;7� �u�=$u	�^�^���Ê�&3���r7��G�=$u���&�����r!
�G�=$u
�t������
��Ţ&����Ê�(3��r7��G�=$u���&����r!
�G�=$u
�t������
��Ţ(�����V�
 � �<$t�FG���� �F��^Ê�` �}$u<0t<1u�`�����6 �Ê�a �}$u<0t<1u�a����Ê� 3���r7��G�=$u���&�����r!
�G�=$u
�t������
��Ţ����Ê�!��}$u<1t<0u�! ����Ê��6 �}$u<0t<1u��6����Ê��6�}$u<2t<1u��6�<0u��6 ����Ê��6 �}$u<0t<1u��6����À>�6tC3Ҋ�"r:����G��r-
�G��r#G�=,uG��������6����6���6� ����<1t<9uH�}$uB$��������E�}$u-$
Ļ�4� :t������GS��6K���6[
�t�2 �����      	�( ���������������S�W�_S3���&�&�O�ډ�O[��&�G��*&�[À>�6 u/3�Ƈ�6������6CƇ�6C�p���6��6��4��������ø@ �l ��&���&�;�t�3�3Ґ&;u��s��� s������ �3 ù	 �������X�Z� ������ZX��������ZXø@ �l ��3�&���&�;�t��&;u� �������X�Z� ���������s���v�ZX�)ZX���6�@ 3����6&�F< t�<
t<t<^t�G&�F< t<
t<t<^u��$��6�S�؀�0��	~��߀���
|��~�����[�S���6�[2��	�!�2���!�SQ� ��P$�'@'�����X��Y[�PSQR� �
2���
�tAP��PZ�ր�0����ZY[X�                         �                                                                                                                                      MITSUMINOFASTDISKNOSELECT�79F:�<�;{>�?@�?�?@)@	819{:2=�;�>.8X9�:^=<�>�8�9!;�=�<B?�8�9J;�=�<b?�8�9U;�=�<o?�8�9w;!>�8�?�8:�;8>�8�?�8:�;�8�<�?�8:�;O>�<�?�8(:�;`>�<�?�86:�;m>�<�?
ATAPI IDE CD-ROM device driver version $WARNING: Invalid parameter ignored: $
ERROR: Unable to detect ATAPI IDE CD-ROM drive
ATAPI IDE CD-ROM device driver not loaded.

$ drive(s) detected
$   unit $
# Monaural Audio Play Mode
$MASTER, $SLAVE , $polling, $I/O address 0x$, LOCK$, UNLOCK$
Driver lecteur ATAPI IDE CD-ROM version $ATTENTION: param�tre invalide ignor�: $
ERREUR: lecteur ATAPI IDE CD-ROM non d�tect�
Driver lecteur ATAPI IDE CD-ROM non charg�.

$ lecteur(s) d�tect�(s)
$   unit� $
# Mode lecture audio mono
$MAITRE , $ESCLAVE, $scrutation, $adresse I/O 0x$, VERROUILLER$, DEVERROUILLER$
ATAPI IDE CD-ROM versi�n excitador de dispositivo $AVISO: Par�metro inv�lido ignorado: $
ERROR: No puede detectar mecanismo de rotaci�n ATAPI IDE CD-ROM
Excitador de despositivo para ATAPI IDE CD-ROM no cargado.

$ Mecanismo(s) de rotati�n detectado(s)
$   Unidad $
# Modo audio-tocador monaural
$MAESTRO, $ESCLAVO, $Determinaci�n, $Direcci�n I/O 0x$, CERRAR$, ABRIR$
ATAPI IDE CD-ROM Ger�tetreiber-Version $WARNUNG: Ung�ltiger Parameter ignoriert: $
FEHLER: Kann ATAPI IDE CD-ROM-Laufwerk nicht erkennen
Ger�tetreiber f�r ATAPI IDE CD-ROM ist nicht geladen.

$ Laufwerk(e) erkannt
$   Einheit $
# Mono Audio-Abspielmodus
$Sendeabruf, $I/O-Adresse 0x$, VERRIEGELN$, ENTRIEGELN$
Versione ATAPI IDE del dispositivo di comando CD-ROM $ATTENZIONE: Parametro non valido ignorato: $
ERRORE: incapace di riconscere il drive CD-ROM ATAPI IDE
non caricato il dispositivo di comando CD-ROM ATAPI IDE.

$ riconoscimento di drive
$   unit� $
# modo mono di riproduzione audio
$ELABORATORE CENTRALE, $ELABORATORE SLAVE   , $indirizzo I/O 0x$, BLOCCAGGIO$, SBLOCCAGGIO$
ATAPI IDE CD-ROM �f�o�C�X �h���C�o �ް�ޮ� $����: �p�����[�^������������܂��� : $
�G���[ : ATAPI IDE CD-ROM �h���C�u ��������܂���
ATAPI IDE CD-ROM �f�o�C�X �h���C�o�͓�������܂���ł���

$ ��̃h���C�u���F������܂���
$   ���j�b�g $
# ���m���� �I�[�f�B�I �Đ� ���[�h
$�}�X�^�[, $�X���[�u, $polling, $I/O �A�h���X 0x$, ���b�N$, �A�����b�N$ 
$IRQ $, $V 1.54 (11/21/1996)
$V 1.54 (21/11/1996)
$V 1.54 (21.11.1996)
$V 1.54 (1996-11-21)
$Copyright (C) MITSUMI ELECTRIC CO.,LTD. 1994,1995,1996
$                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        LN   : F H N   edit.hlp          F   b  �  s     �          �E  �  n  �  �    �    �  g  x  �  v  �  "  d  0  �  �  �   O!  �!  �!  1"  �"  H#  |#  �#  ;$  c$  �%  �&  O(  *  �+  U.  ~1  .3  �4  H6  #7   8  (9  �9  [:  �;  S<  �<  O=  y=  �=  >  5>  �>  �>  ?  �?  �?  @  r@  �@  hA  �A  B  �B  �B  C  �C  WD  �D  /E  �E  -916 h.pg1 -917 -902 -904 -908 -907 -909 -913 -365 m.f m.e m.s m.o m.h -288 -289 -291 -292 -297 -299 -302 -303 -305 -304 -315 -318 -317 -340 -341 -349 -350 -351 -9995 -9992 -9993 -9998 EDIT.COM EDIT .cccp -9994 -2007 -2014 -271 -2025 -2024 -2027 -2051 -2053 -2057 -2061 -2064 -2052 -2068 -2070 -2071 -2072 -2067 -2076 -129 -180 -254 -265 -255 -256 -270 -219 -218 -2075 -245 -215 h.pg$             	 	 	 	 	 
                       ! ! " # , , , - . / 0 1 2 3 4 4 5 6 7 8 9 : ; < = > ? @ A B B C D E E 	$replaces4The5The5Use7The8Each8You999399949The9UseAllowsAltArrowBack	BeginningCancelChange	CharacterCheckChooseClearClick	ClipboardColorsCommandCommandsCompaqCompleteComputerCopy	CopyrightCorporationCtrlCurrentCutDOSDelDeleteDialogDirsDisplayDownDrivesEDITEditorEndEnterErrorEscExitFileFindFoundGettingHLPHelpHomeInsInsertInternationalKeyboardKeysLPT1LastLeftLine	LowercaseMakeMenuMenus	MicrosoftMoveMovementNameNotOnlyOpenOptionsPagePastePathPgDnPgUpPlacePressPrintPrintsRepeatRightSaveScreenScroll	ScrollingSearchSelectSelected	SelectionSetShiftStartedStopsSwitchTabTextTheThenThis
TrademarksUpperUseUsingViewWhatWholeWithWordWordStarYouaboveaccessactionactivateagain	agreementallalreadyalsoandanotheranyareattached
attempting	availablebarbarsbeenbefore	beginningbelowbetweenblankblanksblock	bookmarksboxboxesbuttoncancancelcannotcasechangechangedchanges	character
characterscheckchoosechoseclickclosecolorcolorscolumncombinationscommandcommandscomputer	connectedcontainscontentscontinuecopycopying	copyrightcorrect	correctlycreatecurrentcursordetecteddevicedialog	different	directiondirectories	directorydiscarddiskdisplaydisplaysdocumentdoesdowndriveediteditingeditoreffecteitherendenterenteredentireenvironmenterrorexcludeexecutedexistingexitfilefilenamefilesfindfirstfloppy	followingforfromhardwarehashavehelpherehighlighted	includinginformationinsertintoitemkeykeyboardkeys	keystroke
keystrokeslastleaveleftletterlinelineslistloadloadedlocatedmakematchmatchesmaximummaymemorymenumenusmonitor
monochromemousemovenChangenDevicenDisknDisplaynFindnGettingnHelpnInsert	nKeyboardnOpennOutnPathnPrintnSavenUsingnamenamednevernewnextnotnumberoccurredoneonlineonlyopen	operatingoptionoptionsotheroutpartpastedpathpieceplacepointpointerpositionpossiblepressprevious
previouslyprintprinterprintsprogramspunctuationreadreboot	recognizereduce
registeredrelatedreleaseremainremoverepeatreplacereplacementreturnreviewrightsavesavedsavingscreensearchsearches	searchingsectionseeselectselected	sensitivesetsettingssincesizesoftwarespacesspecialspecificspecification	specifiedstartstartedstartingstillstopstringstringssubdirectorysubjectsuchsupportsure
surroundedsystemsystemstabtargettextthatthethemthenthistimetopictopics	trademark
trademarkstype	unchangeduniqueuntiluseusedusingversionwantwaswhenwherewillwindowwithwithinwithoutwordwordswriteyouyour���� n l &  l�  +� /� ��$ " b��M�F , �8 2 N�6 �K�D > =�B ���>�j L Ād V T ?���^ \ ��~�b ဩ�h 5���s� �v t � �� � � � d�� � � � ܀耐 �����8�� � (�� ��"�� ���� � c�� <�� ۀH�� � � ����� � ��X���� m�T��h��� a� � � 4�C�� D�� }�� �� � ��ƀ���1����������Z�VT&��B@642�����><��Ѐ��%�RH��PN��Ȁ������Zf��xvljh��؀�tr��̀ŀ^�������怈�뀒���ɀÀU��
������r���g������A��Q������р�����Ԁ'�o�: �e����w���\�z�������3�� �*�P�߀����`������#�$n�86,��42׀��R�u��B@i�.�fTNLk�L�R��7�`^\Y�	�I�d;��������t:�|z�&�����ހ������ـ��΀��]����������Ҁ���{��������_���ڀ��π��W�F��j�$�t��H&��,����q���)��0�6� �����J�E�@�Հ[�����$!�S�F@20��6v�><x�V���Dp�������|rd^\��b����lj��Ӏp��݀v�z���������������通�������ˀ���ʀ�������������������̀�|��G���h�B��9�y��-����2��O����  � pO�m��H��f��
F�t8���O�<��HЂ��Һ��q��'�Lf��ϙ����RlZ����)'=t�(��m�~4L�ط�3B/�?�`(.�8P��D��R4 �8#����j��HK9*c48���D� zWF�ڎm\^sZG�2�i ���?�9�~���i���G5�&�r������V���[G�� ݺ:�c�l�G44��-���#����:8e�ѣ��`-x9�	�R���2�(F��Eѿ:؍��� �#��hP����cwH�YB4
(F�����7:>��%��G��=�:�>1��	]��;(� 죘�x�#e�O�ԺYP�S�+��&#t�8G?����c���u�E5t|��6��9	]wu9 ����/��;�@�9� �uɅ'��?ϖ�s�i�����!%H�j���Or`����!��.lo n�t�@C����*c4=�"��v �J���Q�Ӊ�4��9�E�����]lӗ-qS40���D�ĵ �(F�dQ�i�I��r���2���=���4@E�ĵ�g澇�j�r]2�h`�WF���o��p���tw�B4o9��bT~���]]�P��(����1��º�;ҡ7��u��7��+�GG��F�9��;�t��.�BW@��pG�S�Ԟ�7�`�:>CH�)8���j9�bJ9�OY�e6H������t��yut�u���'�%�H��� ߑ���u �+��sy<n���E9Ч)2|d��򜉩D�t�~�T���L�ˏ���"z��ZWH m���Y(��,]dn%� �#��<F�<��+�ts˫�ˬ��46��=�|��9�؍�|��At��@vQ�����oHЂ���h�I��f�G���l�]
pr������&*��T�Ч!���kt�:`��2],|��	b��\��
L��>F��t~bf�t|�=G�	~�MɁfOL|C[���	��G�>�.�>B�����C�~'D���*c1)��(q��j����Q�]�TX�D�9`�b����R��=�;�����8�ʁ�R�=:9`���#p$}I�����9�b7I+�ӣ���#��k�b5.�T%��J뻡��H��إ/�;`X�����0�#f'm{`ڠ;X��%t�a`nD�❰�B�;�X5O���0N?��ށ�K���ibN����x���\��U�+��@����1�:!q��A�I��Һ=j9�q���X�D�9`�b����R��=�;�����8�ʁ�R�=:9`����BH0�P�,��o��N]+�ӣ���.�7GԞ��M�����#q���=:9`��2�J�܂���1�sRT�i��9��Kp��}�c.�.�X:�`<�f7t�sX;v���W]�-H�GԞ�)��X'h���oda���lTk���� l,Ȕ@��S�(X��'u+��0�I�����2#�t+K)��Б]S4���x���\��U�+�S@���e��v��)�,RV~ ����SWG��]  �T�@n���@'F1���?��wB�&�ZWH�����=1^�c1�?�- �=�\p����kJ맳�"� :3�<�&3{��j ��� �<U�+�@C��u�1�Z�2E5����
F�CbWR�m�� �sX��8GX�Qͫ����ë�R:&ES�����lck������kmY��Ԩ9JI$��� e�-�#|���S�u�̜VR��P���B7�:��I$�N��~����h5�1�$��P���B7�:��M]'��ts��s�B7�e�,��TCT��~���
�o���Y�ԩ�::m�ԩ�:�ڎn�G?H���T��F�[a����	5�s����S��7��O|��7A�Bs��1���GGL��:$"g:��-���Ŋ�:tt�=$�c3�ů�-|	2\��bja%�c�뻤 �!1��N��8��c4\|��3G��7�:�@^t�u����g`�,J��M�1���;�.��L�u9��,E*�tf7�yz��h�a&n��L	�+��%�1I��A�M\Nʏ�躚@�L�/�0� +�C�~bi@к$[��R4 �()L|��4@="F&��&>A���՞���_&��w!,B��U�eԪ��?�(�NC���$���3D�>�4�%\�<1k����ɫ�э���H���W	��:�� n�t��j9��NJ���X�Y��ut��9��d��M����c��0�5]"]�u�z����2��Ջ "�a6 �ۣ�h:� = #.����m�d��JW]�d?�Nt��R4 �����= #�73u*t�dO�|L����!� �+�AA�|#B
C`i�#���'rH?u�����1-�w �4�����n�
�cx����f7�x���tg} �A�'rH�1��A��BY,oG��+�{j�W�u���䩌����Y��;�"�⢫��M���L�*%��!��X��;;�)T]~:1������ �+�����W���bq�|��o`lLĮ�;;�)P��OA�]o�A{��3G�� h��wS�	��Ĭ|� �bv���o�4J� �H]=�S��}\F���3D���n������wKY�O�V?ֺ� �bt�� �+��E�NJ��h�;,s�N�W]�"I?HЂ��?�%)@�7:&@��h�z�c�4$�)�}\F���y���߇�W�/�!���ׄz�����>3���m3]T��� @^~ ��E�5f��)�h���ZA�U��]�j�O�=�,K�S�h?6��3&��H-Hm�Pr�&@�\Sd����OKаc�� �+���-#tOS�HuvwĲ��t�l�2��s��8$�+����&Aԝ����oHЂ���h�I��f�G���l�]
pr������&*��T�Ч!���kt�:`��2],|��	b��\��
L��>F��t~bf�t|�=G�	~�MɁfOL|C[���	��G�>�.�>B����aT�p(�J��A��
F����wG�Nt)�hG���,L��ꙃ�v�#B
C����9	]"vw�R���tc��
p��/	]�w�R�l��3{!N��WG�w�R�F1���>A9" A�t���C�N�W@~j�T� QtNXM���/���1�%c��"�j*�fL��t|#����EX��0m����xwҺ��2B�7D���M�_�c������.���t�H�%��C�7�G�Ax���]wu*I��|h[lWG����_A��WE1�3-H���<7���j?G�5�*)��]�W]�#$?��!���I�3G�o�'L1Ώ��@��%�%4���0�h��k���31��~�:`#����"T�`Qt|�#���<>�|u�f'� ��a?u�)bM��֚��A�|a�]wt8!i�}]�Y��/�����y���#3?�Y��-#t�8p�o �]�hAy���u��2A1S�A����Џ���4|��t����D��_�S@Y)]wu*I��|h[lWG����_A��WE1�3-H���<7���j?G�5�*)��]�W@�@�%�
.��K4��<�����G��N/c�!�שN��<�f)�M�� h��wA�b<���Џ��"f����C&3y��yן� �P,�]wt��f��BLs��$�vc�#���83GAJ�+���&*H3
��Պ��G������7&.���鈙#��o ���ym�=Θ �G�5�!31�k�4�J� @�(��p�M����������/���on���&f1�>��&���`$�Cx�Ԯ�� ��]-IS�8R����%�ZF�k��K�f~�x�,u��cy���녁�	ڕ�wC���q��G�@"�� @C���������A�8�'�J뻤X��7O�z��W��,u����녁� q+�������,7��%<|�*|i箕��g|ORzD���o@ni�ׄ�J���RQr{�E��*RQr{ͱ�͋Q�1�:q��\�U��Ey��1��,�����T�Ov7�@"���2�s�f'��!"��4�Q&n�0�#�����%�'�J)�@��z.Z�m������pvwĜ��I��1T���;�N���I�`����)2|*�2�\p����W@� @^~`(�@���ة�������j��i],[;�[d)��������'1Ή�5��~x��e�Ə�L��wA�B�Rxz�D"SW���z.��+0���#@J� @��,M(]P�b<���#�����ND��bSq�HЂ��#��bW@A��S����T�bSq4�I����;�d��R4 �w���!�8P�;���]�����y�0� +�����8��H�R����0�),��1+�� C�~�(�A�1���M�h~����6�z�b����%2)�׌�5t��R4 T��;;�R'�<��5�-���~�����ti @�i���
.�IS�X��t��K+��A�1�H�R�]@C�)6-LZ��qI9��wt���0� �MU�h����G} �Kj?�`)R����+���G} �Kh��  ~���z Y	]4�j;�h��;�@@���)�,����5�3Z�b�W?��9a��������<��J��sQ�H3~�8?@�<R���u�M�o�j������hAJpG'�j��hwu�9���1Ώ��#c���YN�7��q���t�,�9��t����z��1�:��X���L != l�c��U�D�����hAH O�ժ���]}�'H@PN�'8�HЂ���n��L  :h �Xl����׈!Wũ��bj��5 �HЂ�q�T��^Wܒt�
*����LT�|/�����Cp�||��%t�@^~<�>�od!�'��4���*����������R�� �{
*X�CTQϮ�3�h�&a �G�#@J���9��6���O����� �@B`'Z���N�I0�
�g(�sQ	�l � �SR�����8���0Y�TԾ�}�$�C�NGHsQ<#B
� �*���!ܒa2{9�����@>�SR����M ����l �!u7����� � �@����]}��u�}��t)}���y=��,C!�	(��t�Ĭ|�b����+��G��c4#�܂ ����وl `�	p���H�p� z�I+�@u�E�A������Y#�b�G�Å	�/I�����M�6e�8�D|�a��W<�B倲8���A�Ciނ��s@-���	�#�
w�O�x;���$p���zLf ���w^1���/D|��8&'>K �p�����Rl|F�m9jK!���	]wuш�"8P�M8Nz�>Y#�bq �J뻮��LT�.�}�ܮ���_v�f����#��G��R��W��G�c�#��E5 �M\��_y���z�q��a5Z�|Е��B���h�,��@Bz ��@  � sUw�������/� ��R'����d5A%��ؓ�0�)������t��!�t��d���6bh ���𝤒G5K��ԒI]x���
(�PT]1����p�J#���a�\1?t��)MQU#8o���9�W<邓'�M]��p�AA�����u���%thw�;�J뻤V"}\ �:t�b���
Kb> �H�ԡ6���k���a����z�H頃�U�G�����-@�G�>����J뻡�>��H�B�G�pR;�R��WC�$��8r�>Jh%+�AI�s������#s!#�bT��f��H��s�r�#��Lc4|����H㖢}]����\ڕ�wA�D� ��G�ȑ�5��'�X�#����h�^Z���}]���uZ�9u7����� � �@����]}��u�}��t)}���y=��,C!�	(��u�bg���hAA8~뻤Q�G} �ֹ���ϫ�#B
X~ ~cx��9����t�|��WG˖ �czT��!@�c�+�5�0�5����R4 �8#c��ܠ~��'�gL�%�c1t���D1�����t��J뻩Ú��A�.>Rbqt|����<�8J뻠��G} �Ķ����@<����������G} �)1����;��<��ޏ���d1�׃�#�8 �S��/?Ce'������Ÿmw��u�:bm2 $U����sQ�H3���ȃ���I�5��+��;�"���lx�7�lG�5��%u���sQ�H3���8$�~��x�u��;~����j�h��'✆�dZ��u祤��$��'@�z}�9��[�P5z1A:k��a+��@���
F�wS{ != l����T 9�����]�^W�]�B�ܐQxPN���PyR��2���}w^1&C�ڒ�h�Ji�"���Pى�A�HЂ����{�%�ZF�)G�� )�Ϲ1v���<�3�?����'��1�NA� �~뻩�Cƨ���W�4x0��5}e�_^���xj��=wt��16*pL�_�m�*blV��P|�Py{�F �8Po>M�����X�������3�����CG8Ho��a�s�[$EY�f/�ġ�)$I��=Ԡ�[o��ӗƖ�s�ğ�kC�C���R4 ��u�9i��$���pI���ٽC�8A�Ə�
F��e!Y=��=���_���H㖑�mn���hX�O"���j�ƃx�4�$��ȧ8I��-#�¬[��3����G��j��+��Z8����h �Ci�E!Y��S�~	����e׃��8)dS�"���v��_�}\!�~mxE�������{�a����e8@:�G��Ps�q���t)�����z�^���t����?�I�7(y�a���wA����b�𙁄�u
S���I��L`�(�+��=T�SkO�my����p	�dM l��j��U�t.�������䂈uH<�ʖ����s����)PJd_16+�WCh�1��,�S�� ���shymqV��uL��l��L��31]���%���+h G��h�Ķ��^~M]!�Iܩ6�|ן����y����NZ�� �cyV+=>%��<Җ$�`�n�9�<b�����*���,I���-��}Yk���]�3�?u(�Җ$�T��̻x��A��c������-�+t��UI�Vp�	n�hX1ΆGHCR�{��ͮ*�'�K^~cwCf�6��H�a��ɫ�j	L�c{�1�k"���?/���N^czEya��N[�t6�A�����ז�禫X���<co���!��m5ů��Q��c�JJj*�ث8\~�{[���.�]���6+�� 9t.�+�)�`Ă��{H�\�"�����+���!��q���VEuL���ͯ���,�د�n�[M�i���M���1�z�j`�	�!:A8N�
��V�]wt�6�bpH8?<C3����d'J�8&i��@���]�j�Һ���������<#B����%u��۱ 4|�خ1Ə��r:hI�1��ܮ�1�͆���P]�B(5�,˷���4�؍ibN�s��+��h=Ô�ж�cL̟U����3�r��)6���� vз1�>#����{l]"|g�NGs��' +�"�^2|g�NGs��*R�5W���a��_��v��]wt�ؔ��?�r8c��9m�fm��A���ψ7�M쀄8����6@@5P�U�t.���p��t)}�������s뺔bG�ڟz�&֪���5"eWũ��b��	�!O�p�^�4�����h �]wt?�w ��Bx,T��w\��`6�̖�fB 8o@@��@T��KK�����rI�Z4Z�@ pt��:��$I��������]}�}�'B��2�����L #�I��RE� (��zB p*�/�@����o�䓤�h g��L  aH�� 0��� ��������S� Wܒt��=��g��mğ���hADq�ń�/ȧ��o� a�3�u4�ry���A�:������1)w]x�xZX��Ű�#w�}i5t��R4 ����м���?�v[�����\);,�X o����@���%���u7����� � �@����]}��u�}��t)}���y=��,C!�	(��t����Jj���p���`=��Z�hH�brc0?���"�}�u���w�>����vα��8o dx}��XvQ�hx�#�u�4 �^���6��j9�,]#�u���G��X���Y�'�"�� g�J<ٝ]#��s�9�)(
lk�]#�6��/�嘚�j9�,a�G9��t��� ��P8�� �얎�����15Z�sP,]#�u�g���>�h�:İ'`��}����;a�G9��bX�A�c� �pL�m(�_:�Glm�!�'s�c:İ��_�v�]#�u�J�w �4��cc�:ΰ���/����8I�ut���!�'��_�c�:ò�sC�顰죜��bA���e&�caI����� ��6@@t��� �]�B����+���K�H(��('T���(<�`zPIG>���!x�� �`Z� ϱ���!x���"E��9 Ϸ��s�����M0-� ϶��s�� ϲE��8P>͗A�A�!S�A\�ސ�.���@qC����hs�>䫠��}wOlM�ɫ=uL|�خ������� �p�7H�B�9�� >�z ϶�x��s��tz N�����n�X�c� �vG�m(���IG>��V�`�c�$���>�Q�e�+�a���s�����m(�*����h�	58�`�듑J�mw�_B��8��&�zA���}K���z�-���}
c�v����߄�R��C�}P�E���C�O@  :hdU j���u�W}ו�W}Х�$@^�A��T�=��$��]�'iHT� ��
�-	�3��]"q��<�g�,�Z(�o��$�*r�. ϵ2��$9�
a���{]�s����	58@� �׼H� $�� g�ˠ��}wC�y�����Ls�㣅 3�<rkt?�f��~r�>�Q㐫[�C�}P�躛�p	�dM l��j��U�t.�������䂈uH<�ʖ����s���>N %�&��OB�G�/�"�Z]rq �:/�}�LK��#@��>���$��]�����x%�%�K����8�/ۈ+���Y�U!S���b�g�5@�uA/�˯] �F��p'8A/�}�3t��f �1�D�_��W@|A��8H �`躛�p	�dM l��j��U�t.�������䂈uH<�ʖ����s�EbrA�#�A��6�=}"���p��"��,��J9��r��q�Lf����x}���IG>����� Ԃ	�f1�>��/����#�;H �fc��y:`>�{��#ь�F9�H �fc��y8\�m(�^�$��]��ĳG�v1Ώ���x%������ ��} ���L"�w��[��H����-��&g8��}wA%��0���� g��<>�;��cj�T�@躛�p	�dM l��j��U�t.�������䂈uH<�ʖ����s�1���>X�G�&8&W�W�p�}�.��G�@���4|c��v�p�g�r�l�z���f9����'�b��rA%���G��!���� ��D�=}w禫^����<t�����SA��N� �E���C�O@  :hdU j���u�W}ו�W}Х�$@^�A��T�=��$��]���Jl�<?"���}���ŭ�\N1JD58�3�l��AN8>�Q�;�/���XS{ != l����T 9�����]�^W�]�B�ܐQxPN���PyR��2���}wCf!R�b�?�`)Pȱ����%�'�Gr`5����8�pN����}w]�Hp	�`K�lx�"q��8X��r����}wA�R�����w;���_���3@R�w8^	~��u����h���'j�� �����l�()1��� w�8�T�@K� ������!X
S�;��MHW��p����ٱ��ޞ�/?�b�Pw&?*�F�]�s����Ǣt���D� gٱ�t��+��;�����'zA/�}�7@e@�h�;��,l1u�������M�;�&������7�č��6w��D##�s�S�����+�ƛ8��`ئt�WS�
&��;�%�lEE�0)b5�L)������NA����s�����s�T� N��gg|A9B2?1�'o�6�J��8P�c�
pr���>�Cc�_2�<#B
G��T�r���ϙ��R�@���#��vwĜS���%�]+�������t��=9o����k���B�b�],6wĜEX�]���J�k��$�s-�?���p��&��cI�'�g
@�#��	] � @C�) ���M.�I?HЂ�N~��ז�b��<���-����y�Ə�9h6��k�\�ۑMU���X����p��]QNtL������� �~ ��~�n)�ڌf���.��H ����Uۺ+��|h�1�|Uv��7�3'Ƈ��Uy���tm @Cꢕ1v����V��5L]�_�#k�	�������)~}�y��\U����c0�] � @C�Ժ���rQJ��x$Apr虉)���2�nP�O���1�:�����O��������R�|L����F�!̂ 7R�q C�~^�,��$�����,���$A?�rk�pP�.�|A�W@� ����b��t|	��O�Ze�b�Xo6�H�+��%�c4=����4bdI),BK�1�����r���Ф����M���@9	] � @�??�m�vCZ&bJ'xc4�&�R����.W����-ן�W kp�Х B������vKf&_0��EL^~1���|hy����N�C���>KT�bȟ%����],D�F3B��+�� @���.܊|p��U�My�G�j��1yS4r�篌f��1�� x�m�/,������c3�G�XX��J뻤L�3��'?G�{���[s��?@a�G�����1x���ހ����������U���.���
���bW@N @C�0]E1w�.����c��p�7�f)->2j��9�t� C�|I��������O
��'-��?}o���,����$����?u9�`)R7(y��|���s����	����1�@�X������t��Ck�S"��>N�$���� @C��1��M@���bYf1�D��h�=)��N�f �J� ��>-_C[g�ב�?DN��,���H�WCB�4G����,�W@� @C��.�97R�����hAc�)*����3��õ"IWH������)L|�!��x>0	]rK���J~����t~��+�4B��d�)�3H1��mk��
F������xo�V6blW1�~�"B=qg-u��8�`�s�ǓW}uZ��u���T��q����-Nz��4'H�|��~����$@���G��)Ά��\�&�б�����t� ~1��'d �W�15Z� zWo
��b�f9��t� AꄅWm�b�L\wRM���T�G�#ZRr7�3�w��oC����X�$������y�Ə����t�з C�}^�bq�m5Z���C��"9R�"�4,q2M&~�Ov7�@"�b�)6�1�>Or�5�	ːAg�ÌJya�3��kҡ.�BW@'AA�p�S���/�f�"*e����mw+����Ч#Ĥ����Bƙ�Si�>?1�?�cL̟:�3�]wt|��>>M���H��*�o��b�>.�����x��c�WK*�t%�?@it<����.p/)H�)] � @^}_�,7��M�
x
F�[�?C�)��8�II]wtH�I�D�3G��o���0��א�Į�{ @^~�X��P@�P�����Kd���1t�&Rd�����~|�����pG���8@^}W����y����ɴ����Yo�hÁ��%t�؇�~L�O	� �Ğ>Md���0�||�@D%��B��O��0'k��"f���oG�#B
$�,J����:$A����n6�8�E+��@���~z�����d��;4'�)�z���t�<��=a�L�A� ~��bb}��G�w�R���tc�� �~ ������Nt|����N��0���­�DT���t��
5�-_&f k%tg|E+�Όc1��<�%�Nt)�4�F(� ��AȏQ�W����t���#�@4J�3��"� :1����"���c.��)
p�%AA����!fk���'�ɣ�&I�I����#����1y��K4�b�n�b�>�����s�y?�����	��#���wR��#k#t�6K��ޅ�&Ll1�f����+p�r�wK:݊_����q��abE+�� T`Uyi�a�D��B]N����Aܹ���v1��A�5.B�v���X�CP��r E+�c��0m�A�8ɫ��jBW@�������,����k�Z��G�w�R���thX�s�d��>�a��j��L��k�D�))��:>CF+�K�<|��p���W =c�L�ث@��p���'����(�������W���f�!b>AܹA�~�p�-�k���; %t���J��bz�<���	��t2p�@�1��%t                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                :start

c:
dir /s
goto start
h
  msg27 db "Copyright (C) Microsoft Corp. 1986-1993. All rights reserved.",0dh,0ah
        db '$'
;
; msg28 db "Unable to load translated messages",0dh,0ah
  msg28 db "Unable to load translated messages",0dh,0ah
        db '$'
;
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               ���� �L ?XMSXXXX0  }     T                       �            x      ��.� .� �S.� ��G v�O�[����Cu1
�u���<u�� �<u��.�>2 .�I �<	u��.�p� ���.�." ����6q� �����/�f��f�����VWQ��P
�t2����rX3����s���>   uR� Z� �>0  t	X3���3��PXP��% ����X��� �y:�>/  tVWPSQ�@ = Y[X_^u�+ �>/  tPS�B = [Xt
3�3ҳ����� Y_^���6pW˴�P�ô�I���p �>0  tô��+< =@ r�>:  u�- �t)� 3ۀ>-  t�@ ;: s�: �+�3ҋڋ>J ���6 �=&�� ��&�D�  � ��VDISK3���&�f � ��� ��t$� .�>���� ����G� t�0  ��0 À��t
���t
.�. .�: ����`���F�F�Fa.� P�U��F�F�~ ]XXt	�`� �a���=�t.�.& �.�& �  .�>   t.�: �  ���<@u;�t!�>* t���>-  t��;8 r	� �* 2��3����* 
�t�*  � 2��3������>6 t�5 �t�6  � 2�ó�3����>6  t�P �t�6   � 2�ó�3���Q�>+ u%�D �>4  t� �u� �� �D u���4 � 2�Yó�3����Q�>+  t4�>4  t4�D �S �>4 u�t3���u� �v �D u���4 � 2�Yó�3���.�>/  t� ��l��.�>/  t� ���ˀQ.�>1  t� �- �'.��.��%x ���|3���H��@� ��t@2�Y�  P�d�t� �`� u1���d� u(� t#�`�"����Y�'���"� Q3�� �d���Y���X�Q���u���I uD���d�@ u;���`�7 u23�.�2 �I�"����d�  u�� � �a�t�� �a�u��� �3��3�� �d$���= tr���� �
�t���� ��� � �3��= �tr䒨t"�2��$�
�� � �3�� �$:���u� �3��= �t
r
�e�u"�2��e$�
�� � �e3�� �e$:���u� �3�Ë�R��?�Z% ;�u� Ü����u�R� ?�Z�u�
 .� � �`�@ ���6� �6� �� �� u.�> � ?퐐����.�> �� �� 2�� ?�a����u��� u���d� u���d�	 u� �3��3�� �d$������u��� u���d� u���d�	 u� �3��3�� �d$����t����� �d$u������ �d$u� �3�����t��R�)�Z� ����u���  u� u���d� u���`�	 u� �3��3�� �d$���.�E � Ü`P�Ў���.�E ��a� ��.�E Ü��m� �u�2 �>2 v�3�ø �     ��SP3����&� ����&� ��[�X��P�Ý��� �[��U��P��3�����&� ��&� �f���Ft��  �"��9Ft��3����&� ��&� ��NX]ϴ���r@&��&�?PTu3&�Lu,&�G��t$��S�P��L�� �F�X
�t���� ���3��3�S� ���&�>P OLu��&�>�� �u�f$<u�< �� [ø$��r	
�u��u7����r9&�G�u(&��t &��#t&��%t&��	t&��u	3���� �3�Î��������������&;� ��������u&�� $u� �3�Î��������������&;� ��������u&�� $<t� �3�ø����&�> �u,&�
 <+t<*u � ���&�>  T1u&� =60t=20u� �3���� �Q.��&�?ZBu*&�IOu"&�Su&����E �G �� �E r� Y�3�Y�� �3�.�	&�?Buu &�llu&� Su&�.Au&��Vu@�QVW� ��ؾ ��h	� �� t�  _^Y� PHILIPS�� �CSS LABVWQ3��t	.�>p	� �u@Y_^�DELLXBIOS �� ���&�> ��6�	�
 ���������&:uG�����3��0&�}&���=  t�=��t�= u&�� t&�]�E �G � �&����0tǋ؃���������  t�&=������t3��� Q� ��t%���t3���t���u	Y�ٸ ��Y3��Y3��Ë����t� ��؁�^� �;�0C�/<�u�E �G �/�OR�^�EZ��^��/s� �u
����D\�ÊO
�I 3ɊO�1 �O���t�2 �w��u
�>K u�^�O+���> �_�t6�>O u/R��]���
�t��C��>2  t�,���2 ��0���.�Z�S�G=u
�>K u�^��[�e����N� ����4�� ��I[ ��� �[� ��[� �	��� �
��  !�� $�� 'B	� '{	� $c�$ �0�N�3	$I �6�	�� �9�� �<��� �   �� �h�        � �   �  EtV{Q�N�Z� H8NM�A�SRI�CrT�              ��ptlcascade att6300plus ps2 hpvectra acer1100 toshiba wyse tulip zenith at1 at2 at3 philips css fasthp ibm7552 bullmicral dell at �3 5 2 4 6 7 8 9 10 11 12 13 13 12 14 15 16 17 1 �PSQRWVU��> &�]
�t��~���3���  �>  &�E� ]^_ZY[X� W �������p�����p&�&�&��0�!<s�u[�� � C�/<�u��[�� 3�P��X% �= ��[u�� �=�s�H��z���t�O �����l�����t�n^�>J u
�+  �� ��O�s�}���T�Z���>H t
�]�t� ��>0  t�i\�P�<	s
�M��\�A�>Q t��}=@ sd�p&��&��&�?u
&�G&Gu��
���<^�u@�\�g ��]�a �>M t�]�T ��!<u�3�� �> &�E.�& ���, ��^�
 � �����.�>O u�# �	�!�.�>O u� ��!�.�O � �	�!�.�>O u.�>P uR�	�bZ�!.�P�Z��ȹ#_�����������= 
r- 
�pÎ�3���������� ���ON����p  ��3����� �q &��" ��&�D�$ ��WVQS��t� 3���&�B � u&�~ � u&�� u	&�>� �s�>[�m� re�6>�Ȏ�� ��F�� �� �� � �F������  ��� �&�B &�~ &�&�>� �u&���� ��?3ҋڋ>J �<��Z�[Y^_ú[�>H�u3����= �t= �ð%�p�q
�t�t��                    �     �� �                3�S.�<���&�&�Bt[&�W�tS��&�G+�SP�� ������B�D�6>�Ȏ�� ��F�� �D�T� �F�����
�tX[3��B�D� X[&�G  &�G�6>�F������ [�SR�: u,���&�&�Bt &�W�t�L��B��D3ҋڋ>J ��Z[�03COMPAQVWQ.�>:�e� ��Y_^�ZDS CORP ��_= s/�������� �u��p&�>�&��&�=t��
����&�E&�E�>&�E  &�E &�E  &����&��bZ����&�D  &�|
&�D  &�D  &�D �&�D �&� &�D  VW� _^&�|&�D
  &�D�P&�L&�D  &�D  W� ��� ���P� �uh��>� 3ҋڋ>J �����P� 3��&�D  _W&�|
&�D  &�D  &�D�P&�L&� &�D  � VQ�( Y^&�D s&�D��_���p&���&�Ë>� ���s3��RQSV�C r;�h�u6����r.�ú@ �� @3ҋڋ>J �M��6 ���&��& ��&�D�( �^[YZ�S� ��û��&�?EIu&�SAt���[�      ��> &�u�XrKt</u�N�Lr?t�.�6c.�e.�c</t-�	��^�l�.�6c�#rt�</u	N.;6cu�F���>���� �.�g�T� r��r�t�</u�N���r�t�<:t3<=u���r�<0r�<9w�3�,0����r/t-<0r�<9w����������� �}�rt���&� ���.�g�d� s�Q�.�g<t<
t�(���.�? t.8t�����.�W���.�N��.�O �.�O�À<Ou+.�Q �.�@ 6.�B q�.�}  ��=ont	��=oft��.�J��V��3۾}&�=�t/�<Ar<Zw &:u
�tG��CG&�=�t&�= u�G��.�����w	��^�^룁�� v��u�.�p&��.�R�눃�@v�y��
��.�8 .�S��n�.�}  2�=ont
��=oft�O�.�H�N�.�}  2�=oft
��=ont�/�.�K�.�.�}  2�=oft
��=ont��.�L����@s����1�;�s���.�: �����.;6�s�<
t<t< ��.�6���.�>R t��]�4 .�p&���. ��]�  .�>S t��]� .�8 �
��� ��]� ���ù
 3����tR���Z��0����p&��&��3�&�&�G&�G&�G&�G&�G��
��&���    ��&��bZ2�Q� ��Yr{��tv�� tq��Q�؍6�P�r^��P�uW��PtP�6Q�$y<u;�L�\2����������٨�DtH���� 3��uBV�u�� r�>J �k�^���D��u�Y��}�����s�r��p&��&��&�?u&� u&� t��
���?�>N t#��&G&�W &)G&�_ r&�G&Gt�&� t
&�G&�O�&���&��.�>L�r�.�>Ow��\�	�!.�.�&��bZ����	�5 �\ ��2���3����" �<.�>Ow��\�	�!�.�.�&��.�p&�>�&��&�=u&�Q�9 Y&���
���.�p&�>�&��&�=u&�Q� Y&�r��
����&�U&�E�
 ������P��3ҹ0����X�����6�D  6�|
6�D  6�D  6�D26�L6�06�D  PSVW�6�_^[X6�D06�T - �� u��u����&�U&�E�
������P��3ҹ0����X�����6�D
  6�|6�D  6�D  6�Db56�L6�06�D  PSVW����b5��UU��������b5�2�u _^[X6�D06�T - �� u��u���Ë�-4_^[[3�6D6T��&�u&�]�
 �������Ӿ]�
 �¾]� ��P��� XP��������� X$�':'.�F����t.�p&�>�&��&�=t��
��.�0  �&�E &�E  &�E&�E  &�.�>0�.�p.�>0�t&��  �����     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   ������     ��� �   �  ����   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                
HIMEM: DOS XMS Driver, Version 3.10 - 09/30/93
Extended Memory Specification (XMS) Version 3.0
Copyright 1988-1993 Microsoft Corp.
$
Shadow RAM disabled.$
WARNING: Shadow RAM disable not supported on this system.$
WARNING: Shadow RAM is in use and can't be disabled.$
ERROR: HIMEM.SYS requires DOS 3.00 or higher.$
ERROR: An Extended Memory Manager is already installed.$
ERROR: HIMEM.SYS requires an 80x86-based machine.$
ERROR: No available extended memory was found.$
ERROR: Unable to control A20 line.$
ERROR: VDISK memory allocator already installed.$
HIMEM is testing extended memory...$done.
$
ERROR: HIMEM.SYS has detected unreliable XMS memory at address 00000000h.$For more information, type HELP TESTMEM at the command prompt.
To continue starting your computer, press ENTER.

$
       XMS Driver not installed.

$
$ extended memory handles available.$
Minimum HMA size set to $K.$
Installed A20 handler number $.$
Installed external A20 handler.$
WARNING: The High Memory Area is unavailable.
$
WARNING: The A20 Line was already enabled.
$
WARNING: Invalid parameter ignored: $
64K High Memory Area is available.

$This program is the property of Microsoft Corporation.             
  ���  z�  �  �  � �2��>   u�, ˊ- ���U s&��.��t!.�G.�W.�_����
��
��и ˳����3������ s��.� t
.�O� 2�˳����3��PSQR��.;�r%.;�w.+���3ҹ
 ���u.�?u�ZY[X������&� �Āu<QVW��3�3�.��.��.�?u.w.�G;�s��2҃�
��Ǌڋ։�_^Y��[�Āu��QVW3���.��.���u.�?u
.;Ww����u.�?u���� t�� u��
���u2�tA�u9��.�D  � .�D�.�E��.�D+�.�E.�u.�.��ָ 2�_^Y˳����3������QRVW���se��.�| u`.�.�| t3.�.�\��.D.�>�.��.�=u.�U;�t.U;�t��
�� 2�_^ZYˇ�.�T.U.�T.�볳����3����ĀuF�QV�g�s7��.�| u.3�.��.��.�?t@��
��.�T.�|
�t��^Y�ظ �^Y��3�˳�3���Āu��QRVWU����ӳ�s9.�| ��u0.;Twjr� 2�]_^ZY�R��Z�t.�D+�.�T.F.)F��3���.�>�.��.�=t	��
�������.D.�E.�D+�.�E.�.�E .�T�R�Z�t$��.+D.;Fwt
.)F.F�.�F .�T�k��t.�E.D�t.F;�v� ����.�t�t.�F.D.�F .�E.D.�t.�E.�D.�E.�D&�w&�w
&�G  &�G  X.+D���ȁ��% �&�G&�OX���ȁ��% �&�&�OVWR�����Z_^���.�M.�L.�D+�.�Tt.T.�U.�E��.���3���VR�����Z^���t�.�E.�D����&�w&�
3�&�O&�O&�O&�O.�D���ȁ��% �&�&�OVW���p�_^���.�D.�E.�D.�D.�E.�D.�L.�M��]_^YY��.�D.�T�3���.��.��V.�?u.�w;�u���u.w;�u���u��
��^��U���SR3��F��F��F�&��F�&�L�N���A�\�u rb�F�V�^��\
�d r]�F�V��^��n��^�rJ.��= uB�.��= u5�^��t.�O�^��t.�OZ[� �~� tH�^���]ˀ��t������^���V�&�w&�&��t/.�tO.�G� ��+��rD+F�V�r4.�G.�G������^ËǺ ��ƃ� ����v�~���wr߃��vڳ���������·ې                                                                                                                                I�   ��    �  ҥ        3 �    ���   ���  ���   ���       � ��        � � ����F�V�N�v�.���.���.�n�.�6p�������.���tPQR.�6>�.�7.�w.�w.�4.�t.�t.&>�.�� ��.�� ���~� w9N�s�N�U�� �˺3 3��ÿҥ�.�&d�.�f�.�h��؋��3����8��ۋ��.��F EE���Ӌʋ����u�  �����������������u�  ]����)N�t�^� .6��.��� .>n�.�p� �e��^� u�.�>�� t7���.�G.�G.����.�G.�G.�.�>�Z[X.���.���.�n�.�6p�.����.�G.�O.�.�W.�.�GËЋ�3�.��.��.�?u�uF���B.�?u<.�G.G;�r0���.;Gr&.�G.G�.;wv.�w;�s��+�.��u����
��t.�E .�.�u.�U��Ā�WVWfPfQfR�K��f=��  v�����f����  v���fZfYfX�Ƌ�_^��Ā�yVfRf���n��fZ��^��VWQfRfPfS�����su��.�| ur.�.f�| t:.�.f�\f��.fD.�>�.��.�=u.f�Uf;�t .fUf;�t��
��f[fX� 2�fZY_^ˇ�.f�T.fU.f�T.��f[���f[��fX3����Ā�k�QV�����s7��.�| u.3�.��.��.�?t@��
��.�T.�|
�t��^Y�ظ �^Y��3���Ā�YVWfPfSf���K����f[��fX��_^�fVfWf3�f3�f3�.��.��.�?t*.f�.ffOf;�sf��.�?u.f�f�f;�sf�ǃ�
��f�γ�f�t2�f_f^��QVW3���.��.���u.�?u.f;Ww����u.�?u���� t�� u��
���uA�tPf�uG��.f�D    �+fP.f�Df�.f�Ef��.f�Df+�.f�E.�u.�fX.��ָ 2�_^Y˳����3������QV�����s,��3�.��.��.�?t@��
��.f�T.�|�^Y� 2��^Y��3���UfRVW����֋�f�ӳ�sC.�| ��u:.f;T� r� 2�_^fZ]�fR��fZ�t!.f�Df+�.f�T.fF.f)F��3�_^fZ]�Q.�>�.��.�=t
��
��Y����Yf��.fD.f�E.f�Df+�.f�E.�.�E .f�T�fR�fZ�t*f��.f+D.f;Fwt.f)F.fF�.�F .f�T�N��t.f�E.fD�t.fFf;�v� ����.f�t�t.f�F.fD.�F .f�E.fD.f�t.f�E.f�D.�E.�D&�w&�w
&f�G    fX.f+Df��
&f�GfXf��
&f�VWfR�������fZ_^���.�M.�L.f�Df+�.f�Tt.fT.f�U.f�E��.���3�_^fZ]�VR�k����Z^���t�.�E.�D����&�w&�
f3�&f�G&f�G.f�Df��
&f�VW�������_^���.f�D.f�E.f�D.f�D.f�E.f�D.�L.�M��_^fZ��]��.f�D.f�Tf�3���.��.��fV.�?u .f�wf;�u���u.fwf;�u���u��
��f^�        ��   �  ��   ��                          ��   �  ��   �                  �U���fPfQfVfWS3��F��F��F�&f�f�N�f�n��� �� �\�� �� f���^��]
� �� �^�����fVW.��_^= �� 3Ɏ���f������.f�6��&gf�4   .f������f�N�f����gf�g�f���g�g�fX�.f���&gf�4   �.��= u<�^��t.�O�^��t.�O[f_f^fYfX� �~� tH�^���]˳�����t���^���&f�&��t,.�?uG.f�Gf��
f+�r=f;�r0.�G.f�Gf��
f����f��f��f��f�f��f�f=�� v೧���������U��P�� � � � uB��9Fu;�~��t�~ɦu-� .� �"��ʧ �Î�$�"��ا  3��؎�X]�X].�.��f�v�f�~�f�   f;N�vf�N�fQ�6���>�f�F����f���&�e�>�f�F�f���&�e�����fYrf)N����f��fN�fN��2���.��Y���� ���fPfRfV��f����f����3�.��.��.�?u�uT���P.�?uJ.f�G.fGf;�r;f��f�.f;Gr..f�G.fGf�.f;wv.f�wf;�sf��f+�.��u����
��t.�E .�.f�u.f�Uf^fZfX���t@�z��<� �.�>
��� -���  �� ���� ��� ���� ���J ]��9� �#_����� �u3��r� %��+����p;�v���u.�6
����p�p� �p��+�&�p�¾ ���.�
�+���G�����&��&�6�&��+��&�>�� ������6 �|�D�D X� �tA� W &��&+�&
�- �.�ﱸJ3��/.9�w�� �w.�ﱸJ�/���t� ]^_ZY[X�  W� �.�ﱎp�_� �+����������+��/ �p��&��� �> ���6 �|�D���I u��&�^�&�s�@&�Z�H� ��&�t�&�v�Ì�&�֧� ��&��&��ۥ�� &���&������˜X �P��X� ��              �#>�C>�c>�>�>��>��>�?�#?�C?�c?��?��?��?��?�@                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                DEVICE=HIMEM.SYS /testmem:off
FILES=30
BUFFERS=20

DEVICE=cd1.SYS /D:banana

rem DEVICE=cd1.SYS /D:banana /P:1f0,14
rem DEVICE=cd1.SYS /D:banana /P:170,15
rem DEVICE=cd1.SYS /D:banana /P:170,10
rem DEVICE=cd1.SYS /D:banana /P:1e8,12
rem DEVICE=cd1.SYS /D:banana /P:1e8,11
rem DEVICE=cd1.SYS /D:banana /P:168,10
rem DEVICE=cd1.SYS /D:banana /P:168,9

LASTDRIVE=Z
��� !Aa�	���!Aa�����!!#A%a'�)�+�-�/�/3A5a7�9�;�=�?A!CAEaG���K�M�OQ!SAUa                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                @echo off

MSCDEX.EXE  /D:banana /L:R


d��)*�t+rov�+�J"&C�p-?��P:-��=�������B!����/
��q���uC�	<e��F�<�I�� ف�����  K O      B    Y��y��������!9l��������u���+S}��(7����`+p+Y�Y�Y�Y�Y�Y�Y�Y�Z�Z[ > u /t not loaded
  R6001
- null pointer assignment
 ���                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                =
=1
/11/1996)
$V 1.54 (21.11.1996)
$V 1.54 (1996-11-21)
$Copyright (C) MITSUMI ELECTRIC CO.,LTD. 1994,1995,1996
$                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        ���� �'D6DUMCCD001                         �    @           $       B@                             Z *     2   Z         +           (                                                  G         C    $   C      @  B@       K           Z         U                            �LD?�9 B�9:�?[@e@�B�C�C ������:'::?:?�:�:A;<<<�<�<.=�=:?�=�>�@�@[AqA�AB     $       UMCCD001 Found High-Speed CD-ROM Drive
 PRIMARY    SECONDARY  Master  Slave   
 
 
CD-ROM driver not ready.
 (A)bort or (R)etry :  
 
 
LITE-ON IDE CD-ROM device driver version 1.03
 Copyright (C) LITE-ON Technology Corp. 1994-1996. All rights reserved.
 
Device Driver Name =  

 IDE CD-ROM device driver installed.
 
No IDE CD-ROM found.
 Please check cable or power cord.
 
IDE CD-ROM device driver NOT installed.

                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        U��.�6" .�6  � P�&��.�6& .�6$ �v P�}&��.�6* .�6( �w P�i&��]�U��5�!.�" .�  �v5�!.�& .�$ �w5�!.�* .�( ����v%�!���  �w%�!�����%�!�]�`��.�>. ~.�.�.�  a�`��.�>0u.�2 � �� � ���.�$ a�`��.�>0u.�2 � �� � ���.�( a��2  �F�Ph< � �Z%�FΌ����F�P�Y�u3����F� ��F�� �V�؊�V�� V�ڈ�F��F�:Fr۸ �����,  �F�PhH � ��$�F������F�P�Y�u3����F� ��F�� �V�؊�V�� V�ڈ�F��~�rݸ �����  �F�PhT � �$�F�P�Y�t� ���3�����U����! �4�� �5�4�6�&4�?�! �4 �5��]�U����6�4�! �4 �5��]�U��H�)�<�(�H�)]��
  �F�������  ������  ��������#���V��F��f�F�&��f�F�&�G�f�F�&�G�f�F�&�G�f&�G��>:  u�� ������U#���V��F��F��F��V��F���W#% ��F����+F�@�F��F�;
sx�F� �F�  �F���V��F��#�V��F��f&�G �f�F�&�G�f�F�&�G	�f�F�&�G
�f�F�&�G�f&�G��f&�G��f&�G �f&�G��:  �f�F�&�G�f�F�&�G�f&�G �b�~�^��Z���V�����U��^�8�G�:�G���G�<�G�>�G�@�G�B�G�D�G�F�G�H�>	 u�� �>8�uj�L�J�P�N�L�J �� �T�R�L�J �� �d�b�L�J �� �`�^�L�J �� �\�Z�L�J �n�L�J �� �P�N�L�J
 �� �T�R�L�J �� �d�b�L�J �� �`�^�L�J �� �\�Z�L�J �� �X�V]�U���2  ��&� �.� �-�H�)�<�(�)�u�(� % = t�)�u��>. ũ>. u�� �61 �OY�>
 u�> t������� ����� �h� �61 j j j j �}���.2 �61 �Y��H�)�)� % = u��>. u�>. u�f�v�Y�>	 u\�.� �#�>8pu�� �	�	�
�t��	$�� ���>. t�>2 u
��&�?�u���&� �2  �>. u3�]ø ]�]�U���.2 �5�H�)�<�(�H�)�)�u�(� % = t�)�u��>. uĀ>1  u�D����D���F���.[ ��H�)�)� %� =� t��>. u�>. t� ]��3�]�]��  VW�F� W�>��������؎��� �@� �F��B� �F��F���F�����u	_3��� �`�� rR���t�F����F� ��3��v��F��N��8�m�F�  �������؎��� �N��8�m�F��F�H;F�w���΋8�m���>��.�#�>8pu�� �	�	�
�t��	$�� ���>. t�>2 u
��&�?�u���&� �2  �>. u�F�  _�F�� _^��U��W����f�>�X�> ���>: u�
��:  ����+ @���f�h  ��� � �j�l  ���n�p  �r �t  WRP�  �>�����Ks�����XZ__]�U��W�T�RV�F�D��F��  ���D��  ���X  �V �����\�Z���^WRP�< �>R����Ks�����XZ__]��  VW�����@ ��{ ��&� u��F� �9�F�� ����Ǉ�  Ǉ�  �F�� ����Ǉ�  �F�� ����Ǉ�  �F��~�r����F� �F� �� �F�� ���؋�x��v�^�� ���������F�� ���؋�v� ���+ @���F�� ����9�zvz�F�� ���؉���F��F�� ���؋�z+ǊV�� ���ډ���F�� ���؋�x��v�^�� ���z�|���  �F�� ��������������F�� ���؋�z�V�� ���ډ���F��F��F�� ;ts�	��N��F�� ���؁�� ��>` u���b�b�^�c�Z�d�V�e�N� �D�u	�R�&��R�F�R��(�}��N� �D�u	�R�&��R�F�R�N�	�N�_^���  W�F����.�#�>8pu�� �	�	�
�t��	$�� ���>. t�>2 u
��&�?�u���&� �2  �N� �R�f���&� tWRP����>��  �Ks�� �����XZ_�>. u3��� � _���  VW� V�6���@� �F��B� �F��F���F���F��~� u^3��s�	�8�N��o���6��.�#�>8pu�� �	�	�
�t��	$�� ���>. t�>2 u
��&�?�u���&� �2  �>. u3�^��� _^���"  �F���F�Ph` � ���F�����F�P�
Y�u�6�F�$�b�F��c�~� u�~�u�G�~� u�~�u�G�~� u�~�u�G �~� u�~� u�G �~�(u�d �l  �f  �h �~�u$�~� u�~� u�d �l �f  �h  �~�u�~�:u�d �l �f  �h  �~�u�~�0u�~�u�f �l  �h �~�u�~�Ru�~�u�l  �j �h �F��F��>dt�>h u�G �F� % = u
�~�:t���ÊF������>  �F�Phl � ��FΌ����F�P�Y�u� �ÊFТ9 �~�	v�~Аu�l  �h �~�pu�l  �f  �h  �~�qu�d �l �f  �h  �~�ru�l  �f  �h �F�u�F�t�v �F�t�p �F�u�F�t�x �F�t�j �F�u�F�t�r �t ������>  �F�Phx � ��FΌ����F�P�Y�u� �ÊFТ9 �~�	v�~Аu�l  �h �~�pu�l  �f  �h  �~�qu�d �l �f  �h  �~�ru�l  �f  �h ������  �F�Ph� � ���v�v�
���V�F�F�F��F�F��F�F��F�P��Y�u3��ø �����  �F�Ph� � ��>f u���u�_�)� % = u���~
 u�~u�^�\�V
�F�v
�v�
���V��F��F��F�F��F�F��F�F��F��F� �F�F��F�F��~u�F� �F���Fi�0	�
��
 �F����V�F�����: ��% = u� �F�P�Y�u����F�P�Y�u3��ø �����  �F�Ph� � �3��h�f�F�P��Y�u3��ø �����  �F�Ph� � �x3��h�f�F�P�Y�u3���� �Q��F��~�(t�~��t� �����  �F�Ph� � �2�F�P�TY�u3��ø �����  �F�Ph� � ��F�P�*Y�u3��ø �����  �F�Ph� � ���F�F��F�F��F�F��F
�F��F	�F��F�F��F�P��Y�u3��ø �����  VW�F�Ph� � ���u�^  �\�>�)� % = u�^�������F�P�Y�u� �f ��� ����� F����E���F3��?���� �����������}���������|���������{���������zG�F�- ��;�w�����u����J����I����-�F��������F�P��Y�u3��1���J���I���H�K �6J�6H����Z�X� � _^��U��VW�v�~�>f u%���u��)� % = u�6��>f u3��N�F� ���؊�x�D�F� ���؊�w�D�F� ���؊�v��D �F� ���؊�y���� � _^]��  �F�Ph� � ���^  �\�F�����F�P��Y�u3��ÊF�:F�t0�_ �F�^�F�]�F�\j j�6^�6\����^�\� �����*  �F�Ph� � �X�F�����F�P�pY�u3��ËFFth�F����^&��v��Y�^&�G�^�F�&�G�^�F�&�G�^�F�&�G�^�F�&�G�^&�G �^�F�&�G�^�F�&�G�^�F�&�G	�~� t�F�R�F�Q�F���F�R�F�Q�F�P�~�u�G��>Gu�~�t�~� t�G � �����  �F�Ph� � �f�F�P�Y�u��>Gu%j j ������u3����G�R�P�N�Lj
�mY� ����U��~sh��hp�j�Y�F� � ����u�D����1  �0 ��D����1 �0  ]�U��VW�F:'r3��e�F:4 tW�F� ����5 ��YVW�؎��D�4 � i�����������F� i����D�������_^�F�4 � � _^]��  3�3ңV�T�R�P�N�L�J�H�Z�X�¢G�F�E�D�d 3��l�h�fh��PY����S�����F��~�(t�~�)t�~��t��>�� ����U���]��  V�
�H�)�>)�u�>1  u�D����D����Z�)� %� = uM�@� �F��B� �F��F���F���F��~� u�� ��������H�)�)� %� = t��v���Y�u�� �.� �H�)�<�(�)� %� =� u�x�)� %� = u �(� % = u�6.�h��u�x�6.�K�)� %� = u�(u�6.���u�Q�6.�$�)� %� =@ u�(� % = t�(u���> u
�>. t�X��>. u��)� % = u3��� � ^��U��V�
 �H�)�>)�u�>1  u�D����D�������v���Y�u�� �.� �<�(�H�)�> t!�)� %� =� u�6.���u� �6.�Q�)� %� = u�(u�6.���u�c�6.�*�)� %� =@ u�(� % = t�(u	���� ���> u
�>. t�f��>. u��> u��)� % = u3��� � ^]�U��N�:�F�<�F�@�F�B�F
���t$���t��� � ����u�D����D�����D���F�F�]�U��V�v��8�D�8�D�8�D�8�D�8�D
�8�^]�U��N���t$���t��� � ����u�D����D�����D���]�U��F�
���]�]�U��F��$���
]�]�U��^�F�<�� ��� �K �� ؀� �� -� �� s1�1�]�]�U��F�V� � �� ����K���]�]�U��F�V<Ks��<s��Ps	
�u= s3�]��� ]�]�U��FF<Kr,K��ff	��<r��<��VV
� ]�]�U��`�F����ʋд��a]�U�� ]�]�U�� ]�]�U�� ]�]�U���^&�O&�  � ]�]�U���^&�?v��]�j j ������u��]��^&�?u�^�R�P��6R�6P������^&�W&�G� ]�]��&  �F�Ph� ��F�����F�P�Y�u�����F� ��F�� �V�؊�V�� �^�&��F��~�rܸ �����"  �F��v��F�P�7���u�����^�F�&��F� �F��!�F�� �V�؊�V�� �^�&��F��F��F�:F�r׸ ����U���^&����
�tx�>h u�^&� �^&��>l t�^&���>j u�^&��>p t�^&��>r u�>t t�^&� �>v t�^&� �>x t�^&� �-�^&� �^&��^&��l �h  �f  ��]��^&�G  � ]�]�U���^&�
�u�^&�G ���u�^&�G0	���]ø ]�]�U���J�j j ������u�d �>f u��>f u��]��6J�6H�����^&�W&�� ]�]�U���^&��N�H�)�)� % = u���>d t�^&���d  �>l t�d � ]�]�U��>l t��>h t�>f u	����u����]��^�E&��^�F&�G�^�J�H&�W&�G� ]�]��  �>l t���Ã>h tY�^&��F��F�:Er	�F�:Fv���ÍF�P�F�P�v�����u�"�^�V��F�&�W&�G�^�F�&�G� ���������U��>l t� �>h t�v�v�j����u�� ]����]�]�U���]�]��"  �F�P��Y�u�����F�u�����^�F�&��F�	�F��s�F� �F�� �V�؊ЈF��F����F��~�t2�F�� �V�؊ЊV�� �^�Ӌڈ�F�� �V�؊
F��F��F�� �^؊F�&��F��F��F��~�v��^�F�&�G�^�F�&�G	� ����U��j j �x���u�d �>f u�)�>f u��]�3��>Gu� �^&��>G t&�^�N�L&�W&�G�^�V�T&�W&�G��^&�G  &�G  �^&�G  &�G  � ]�]�U���]�]��  �^&�G �^&�G  �^&�G  &�G  �^&�W&�G�V��F��^�&�?v���ËF�@�v�P�^�&�� �����\�������  V�^&�w�u�v�v� ��� �^&�G�F��^&�G�F��~�v��~�v���l�>h u�R�^&�W&�G�V��F��~� u�v��v��N����V��F��v�V�v��v��^&�w&�w����u�L�>d t�������� � ^��U�� ]�]��  �^&�v�����^&�W&�G�V��F��^&� u�v��v�������V��F��v��v������u���ø ����U��>j t��]�j j �T���>Gu�G����u��]ø ]�]�U���^&�?v��]��^&�? t&�>h u��]Ã>j t�,�&��u��j ��>j u��6��u��]��j  � ]�]�U������u��]ø ]�]��$  �F�Ph� ��F�Ph � ��9 �F��^&� t�F���F� �^&�G�F��^&� t�F���F� �^&�G�F�F܌����F�P���Y�u���ø ����U�� ]�]�U��>h t�����u��]ø ]�]��  �^&�G �^&�G  �^&�G  &�G  �^&�W&�G�V��F��^�&�?v���ËF�@�v�P�^�&�� �����|�������  �^&�W&�G�V��F�F�F�u��^&�v�����^&�W&�G�V��F��^&� uC�V��F�;Z|u;Xr� �V��F�F�V�- �� �V��F��v��v��_����V��F��F�v��v��l����u�H�V��F�;J|
u;Hr�2�v��v������F�V�- �� �V��F��V��F�;Z|u;Xr�����v��v������RP�v��v�� ���u�����G�V��F��N�L�v��v������V�T� ����U��>G u� ��>Gu�G ����=��u��]ø ]�]�U��>Gt�$�6V�6T�6N�6L����u��]��G� ]�]�U��.�@.�B]�U��`.�&>.�<����м@�������@&�G�:�Pu���>|��0 �>� t�܃>|� �>� t�@&�GP��Y�tg�>� tH�>h u�)܋H�)�)t������ �>(tЀ>�tɃ>d t
�>f u����6B�6@����8���:�� ��:��>Gu�: �@�:&�G�0  ����.�<.�&>�a�]�[S��s�������ـ����ˀ��3����[S��s�������ـ����ˀ��3����U��VW�v�~������_^]� U��VW�5�F�!���_^]�U��VW�%�F�V�!_^]�U��]�U��V��!]�U��V�v��tPP���YX<
u�j���Y��^]�U��V�v� ��Q����$<
r7�0P��YY��^]�U��V�v��$�<
r7�0P��Y^]�U�� �
�t� ]��	�Ĵ  ]�]�U��VWVW�؎��D�F� i�����������_^_^]�� W�����V��F�W�~��������؎��� �.2 �5�H�)�<�(�H�)�)�u�(� % = t�)�u��>. uă>. u�� �61 ���Y�:� �<� �>� �@���B���F����.2 ��H�)�)� % = u��>. u�>. u�b�@� �F��B� �F��F���F����F�  �F��F�F�u�1�N��8�m��W�t�>	 t�-7�
 ���5�
__���  �F�P�Y�u���F� �~�Lu�~�Tu�~�Nuh���F�P���Y���  V�' �4  �F� �3��~�sh��h���Y�F�� � ����uh��h���Y�v���Yj�v�j j j j �����. � �>. u��.��H�)�)�u��)t��>. uߋ:�F��~�tm�~��tg�@�<t	�@�
�uH�B�<�t	�B�
�u6��5��<�t)�'� �V��؈�5 �'�4 ������6'�e�Y�'� �uh����Y�h����Y�F��~�s���^��U������'� ]�]�U��V����t�Jh���Yh��Y� �����=R t��rt
��At��au�V�`�Yh�e�Y��At��au3�����t� �	h�D�Y�^]��  VW�	 �^&�?t	�^&�?
u�l�^�F&�?/t�\�^&�?Dt�^&�?dt�H�F�^&�?Mt�^&�?mt�1�F�^&�?At�^&�?at��F�^&�< t<t<
u�	뀀>	 u�� ���0����  �
�t���p����  �
�t�	 � �	��  �����J�	��" ��L�h�fj�h��  ���f��  ���F� ���u����� �F��~�r䡊���h�f������m��������������~�_^���  �^&�?t	�^&�?
u�)�^�F&�?/t��^&�?Dt��F�^&�?:u����^�F&�?:t� � �G�^&�? t$�^&�?t�^&�?
t�^&�?t	�^&�?	u���� �V���^&��؈�F����r����� �V��� ����r� �1��� �V�؊�Ѷ �ڈ�
 ��� �V�؊�Ѷ V�ڈ����r����2  �F�Ph�� ���FΌ����F�P�Y�u3����F� ��F�� �V�؊�V�� V�ڈ�F��~�rݸ �����  �F� �F� �P�v��N�Y3�3ңV�T�R�P�N�L�J�H�¢G�F�E�D�d �f  �h �l  �F��F�:'r��F������  V�F�Ph��	 ��h��YhM���Y�^&�w&�w�����^���@ ��� � ��0��u� �F�P�^&�w&�w�����h���Y�F�P��Yh���Y3��;��5 �%�Y���3ވF��~��u	���$ވF���ވF��~�)t�~�(t�~��t�F�'� ;�����h��S�Y�^&�G �^&�G �^&�_&�G�E�'� �:h��'�Yh�� �Yh��Y�^&�G �^&�G �^&�_&�G  �  �(��FӺ��� � � ^��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      MZ �   �
��G�                                          ��ENU �NSED  
  �������   � $ G v � � � 	 B
 g � � �   < ^ � � � � � �  - G e p y � �  �! �" �# $ "% n& �' �( �P X	Q Z	Z _	[ c	\ i	] n	^ t	_ z	d 	e �	f �	g �	h �	i �	j �	x 
� U
� �
y �
z  { ~ L� �� �� � !� N� r� �� �� �� � /� @� _� q� �� �� �� �� � J� ]� �� �� �� �� � � ,� G� [� d� �� �� �� �� � � � � � � !� $� &� ,� /� <� @� G� J� Y� h� w� �� �� �� �� �� �� � � � %� /� 9� C� M� Waow�,�-�.�/�0�1�23b4�5�67&8l9�^�_�h�i�r|w�|������������2�8�E�F�^�k�l�m�n�w��������������������������&'( )!*"++,,-;.</M0[1i2j3k4lXmYvZ�[�\�]�^�_�`�a�b�����������������������������+�,�N�Y�Z�[ \!f"s#t$�%�&�'�(�)�*�+����Extended Error %1Parse Error %1 (Edit was unable to access the file
'%P' &Edit was unable to find the path
'%P' 2Edit was unable to create or access the file
'%P' #The system is out of file handles! *Disk full error while accessing file
'%P' -Timeout error while trying to lock file
'%P' 4The drive is write-protected - cannot write to
'%P' -The drive doesn't exist - cannot access
'%P' (The drive is empty - cannot access
'%P' )CRC data error while accessing file
'%P' %Seek error while accessing file
'%P' ,Unknown media in drive - cannot access
'%P' 1Sector-not-found error while accessing file
'%P' Printer error on '%P' &Write error while accessing file
'%P' %Read error while accessing file
'%P' (General error while accessing file
'%P' 1Unknown error while accessing file
'%P'
Error %s Out of near memory! Out of far memory!   Edit requires DOS 3.1 or later. '   Edit was unable to find a match.        No more matches found.           Change complete.       !    Can't backup any further.    errBAD_BUFFER errBAD_LINE errNO_MORE_LINES errBAD_PAGE <Edit was unable to read in a virtual page
from XMS or disk. errLINE_FULL errXMS -You can load no more than 9 files at a time. $You cannot modify a read-only file. OThe file has too many lines.  You can
have no more than 64000 lines in a file.  You must select a region first.  mThere are too many files in this directory.  Edit will
display as many files as available memory will allow. hThis file is too large for Edit to completely load,
but you will be able to view the first 64000 lines. Edit ERROR:    OK   	  &Yes     &No   	 &Retry  	 Cancel   &Help  
 Enter=OK  F1=Help  Enter=OK  Enter=OK  Esc=Cancel  F1=Help  Enter=OK  Esc=Cancel  Enter=Retry  Esc=Cancel " F1=Help  Enter=Retry  Esc=Cancel  Enter=Yes  Esc=Cancel J F1=Help                                             �  Line:%u    Col:%u K F1=Help                                    �  Line:%u   Col:%u   Value:%u J^Q: F=Find  A=Replace  Y=Delete to end   F1=Help     �  Line:%u    Col:%u  Loading %.50P - %u%% complete  Saving %.50P - %u%% complete 4 F1=Help  Enter=Execute  Esc=Cancel  Tab=Next Field J Searching - press Esc to cancel                     � Searching line: %u < Enter=Cancel  Down=Next topic line  Up=Previous topic line > Use arrow keys to resize window  -  Enter=Accept  Esc=Cancel  Move mouse to resize window 0 Drag down the titlebar to open a second window ' Release the mouse to close top window * Release the mouse to close bottom window # Waiting for printer to respond... I Printing - press Esc to cancel                      � Printing line: %u  Creates a new file " Loads an existing file from disk  Saves current file " Saves current file with new name  Closes current file ) Prints currently loaded file to printer  Exits the editor / Deletes selected text and copies it to buffer   Copies selected text to buffer - Inserts buffer contents at current location 4 Deletes selected text without copying it to buffer  Finds specified text < Finds next occurrence of text specified in previous search " Finds and changes specified text  Opens a second edit window  Resizes the edit windows  Closes the second edit window  Selects a file to view  Changes editor settings  Changes editor screen colors  Help on Edit commands  About Edit ! Commands for manipulating files  Commands for editing files + Commands for searching and replacing text   List of currently-loaded files % Commands for setting editor options  Help on Edit &File &Edit &Search &View 	&Options &Help &New 	&Open... &Save Save &As...     &Close 
&Print... E&xit Cu&t       Ctrl+X &Copy      Ctrl+C &Paste     Ctrl+V Cl&ear     Del &Find...                Repeat &Last Find    F3 &Replace...             &Split Window  %s Ctrl+F6 S&ize Window   %s Ctrl+F8 &Close Window  %s Ctrl+F4 &1 %s  Alt+1 &2 %s  Alt+2 &3 %s  Alt+3 &4 %s  Alt+4 &5 %s  Alt+5 &6 %s  Alt+6 &7 %s  Alt+7 &8 %s  Alt+8 &9 %s  Alt+9 &Settings...     &Colors... &Commands... 
&About...   EMS-DOS Editor   Version 0.9.019   Copyright (c) Microsoft Corp 1994.   1EDIT [/B] [/H] [/R] [/S] [/<nnn>] [/?] [file(s)]   %  /B       - Forces monochrome mode. N  /H       - Displays the maximum number of lines possible for your hardware. -  /R       - Load file(s) in read-only mode. 0  /S       - Forces the use of short filenames. K  /<nnn>   - Load binary file(s), wrapping lines to <nnn> characters wide. (  /?       - Displays this help screen. I  [file]   - Specifies initial files(s) to load.  Wildcards and multiple %             filespecs can be given.  About Edit HMS-DOS Editor
Version 0.9.019
    Copyright (c) Microsoft Corp 1994.    No Help � Edit was unable to find this help topic.  Make sure 
 that the helpfile EDIT.HLP is in the same directory
 as the editor, and that it hasn't been modified.     [-%c-]  (R) UNTITLED%u 
Save File 4The file
'%P'
has not been saved yet.  Save it now? Invalid Tab Spacing 5The tab distance must be between 1 and 60 characters Replace existing file? You must specify a filename 	�2
Find 
Fi&nd What: !Match &Whole Word Only Match &Case 	%	�:Replace 
Fi&nd What: &Re&place With: &Match &Whole Word Only Match &Case 	 &Replace 	 Replace &All "	/		 -Replace Replace this occurence?  &Replace 	 &Skip  	�1Open 
File &Name: "-&Files: &Directories: 
Open &Read-only Open &Binary Line &Width: '	%	�1Save As 
File &Name: "-Existing &Files: &Directories: 	%	�HC 	
�)
Print Print to the printer on %s 	&Selected Text Only 	&Complete Document 			�>Colors &Item: 	&Foreground: 	/&Background: .	%  Choose the colors for the item   &Default 	!1	�-
Settings 
&Tab Stops: &Printer Port: 	LPT1 	LPT2 	LPT3 	COM1 	COM2 	!	cBlack,Blue,Green,Cyan,Red,Magenta,Brown,White,Gray,BrBlue,BrGreen,BrCyan,BrRed,Pink,Yellow,BrWhite �Normal Text,Selected Text,Window Border,Menubar,Status Line,Keyboard Accelerators,Disabled Items,Dialogs,Dialog Titlebar,Dialog Buttons,Dialog Scrollbars                                U��VW�~ t%h�+�D���u� � ������£��x���
�,� H�!s� �r����������3���3���������G�G�G���G��G�G�G�G���Ў���u"��������|��� ����Ou�3�_^�� ���K����؋֎��Gt<�G6;�t$�w�D���G�D6�6��w�D�G�\���\�G���Ў�3�ÌЎ�S�[3҃� u�֎���������&�G
�t��&�G�U��V������� �Dt�����Ў��M�D �D�~ t4�Ў������u	��u,������D�\�G�D�w�؉w�Ў؋�������^�� U��V���v��&�T&���t*��t�9 ���  �Ў����t���t�U&�D ^�� �D�\�G�؋D�GÃ>�  u�Tû��?�t������� �U��V�!�Ѓ��u�T �uM����^&�O&�3���tP�-�u&X����tP���uX���^&�G&�73��[P����X^��V���6�&�| t&�t���u��w����tP&�3��
��tI��X����^���tP&�3����	t*��X�^�>� }2���?�u���������� 3�����؈TX������Ў�3��� ^û��� H�!�� |�� �S� H�!r�X��	�3�ø �û�F�����t���+����F�á��ø C�/<�u�C�/�����63�ø �V��> t�� 
������^�P� 2����|Z;�~�Ѓ��R� 	��t��Y��X�À>7 uE�>�}8�>}1� ��r)�������O�����=�~������7�û;G|+G����� ����>6 t��M�� ���u��s��6 ���û�M� �6�V����\�T� �D  �D
  ���\�D�T� ���  u�! ��^�V����\�T� �D  �D  �Z��\
�D�T� ���  u�! ��^��t�Ӱ�8uC�����Ê3ɨt���������+������Ê���؀����� � h��

���uh���	���th�Ph�܅�t�j h���u3�ø Ã>: uB�8�� =�}4�9 r/�<�� ;�r#�>8 u� Z3ɺ��!����r
���8 ���: �û����߀�@� 6�!�������t���� ;�s���������Ã>8 t��� >�!��� A�!�����8  ��G�8������u�F�s���ûG�����6�����>h��6�RSh h  � ��ʋЋ�� B�!� ����r�i�����>����6�����>h��6�RSh � ��ʋЋ�� B�!� ����r�w����
�>���U��>>}�~t� �� 3���  �0�!<s3�P˿��6 +��� r� ��ׁ�NW�s�j3�P����L�!6����6���Ʊ��H6�D�F6����6�g���P6�g
��P6�g6�g6�&@��6 ��+��۴J�!6������PW+�3����������Q3��P �6��6��6��gP��.��ظ �B�P.��ۚ�  ��G�>���uXP���� P�B�� 5�!�n�p� %���!�>� t1������&�6, ����3���s�y����� ����&�, �>��3�&�= t4� �`�t��3��u!��������,Ar����,Ar
ª��� ����� D�!r
�t���@Ky羮���� ����� ����� �U��3��U�� �U��VW� �U��VW��.�Q
�u'��@��@�t ��@��@�z �����b �>���u�������M �����S � �tX
�Pu�~ u�F� � X
�u�F�L�!_^]Ë��� ���n� %�!�;�s
OO��������;�s���Et����� U��� P��>� t���� P�w��]ø ��Y��+�r
;�r����Q3���� V3��B 2���2�����Ut��� P�8� ^Ï���� <t)��&�, ��3��� �3��u�GG�>������ыѿ �� ���< t�<	t�<to
�tkGN�< t�<	t�<t\
�tX<"t$<\tB��3�A�<\t�<"t��Ӌ���Ѩu��N�<t+
�t'<"t�<\tB��3�A�<\t�<"t��ۋ���Ѩu���>��G���B���+�ģ����6�?CC�6���
�u�6���� �3���< t�<	t�<t|
�tx6�?CCN�< t�<	t�<tb
�t^<"t'<\t���3�A�<\t�<"t�\��Ѱ\���s�"���N�<t.
�t*<"t�<\t���3�A�<\t�<"t�\��ٰ\���s��"���3���  �&�U����&�, ��3�3�3�����t&�>   t�F�u���@$�F����	 � P��� ���ϋ�3�_I�&�6;`uQVW�`� �_^Yt&�?CC��
�u���&�]� U��VW�V���;�t@�t�3��������_^��]� U��W�v����t ���3�������I� �>���u���@�!_��]� SQ� ��QP��[��Y���t[Ë��N� r3���]�s�P� X2��]�s� ������]�2�� â�
�u"�>�r<"s< r��<v���ט�|Ê��� � Y��;�s+�����3���QW�Gtc�� ����t+�IAA�w�tL�s	3�����0�?&��=  t� �;�r��u��"��r���H���s3���#�R�. Zs���t� ������+W�G��w
J�B�����w
_YË��GtJ�wN;�v9W�s6BSQ�ގƱ��u� �Gt
Ƌ�+ÎËشJ�!Y[r���GtJ�W�����W�w;w
u�w����t��$����OO��_� U��׋ތ؎��~3�����u��~������+����F�� t�I�������]� U��׋ދv���؎�3������ы~�Ǩt�I�������]�U��׌؎��~3�������I���]� U��WV�~�v�ߋN��
�t���2���^_��]�U��WV�N�&�ً~��3����ˋ��v�D�3�:E�wtII�ы�^_��]��  U��WV�v3��3۬< t�<	t�P<-t<+u�<9w,0r���ҋˋ�����������؃� ��X<-�u�؃� ��^_]�U��F-  �ÐU��^���t�G������U��WV�6��tE�~ t?�v��������-�4�����;�v��9=uW�vS�����u��@�����< u�3�^_��U��W�~��3������ъF���t3���E�_��]� U��W�~3�������O�F��t3���E�_��]�U��� VW�v�Ў�� 3��~��
�t���Ȱ������C���v���C�%� t���Ȱ������"C�t�_^��]�U��� VW�v�Ў�� 3��~��
�t���Ȱ������C���v���C�%� t���Ȱ������"C�u�_^��]�U��3��N��ߌ؎��~�F�  u�E���]�U��׋ތ؎��v�~�ǋN�*;�v���;�s����NO�����Ǩt�I�������]�U��׋ތ؎��v�~�ǋN��t�I�������]�U��׌؎��~�ߋN��F���� t�I�������]� U��VW�~ t �N�It�v��VvV�V
�����x��_^��]ËFH3������ٸ ��r����;�rU���FH�fFP�v�]�ȸ�������;�s��v ;vr������V�V�6U�v�R6u;vt�v V6�U���t�v���ZV��6+uV�v 6�U���t�v���;v u��^;�v6�E���T ���V��v��6�E���΋v �< ����v+v�v +v�r�N �F��F �F��F��N��O��N�F��F�F��F��N��:����� t	K� �� t��� �� u�ô�!� @�U��VJ��!��!@:F���u@]� U��^�H�!��r�ȋ^���2��������� U����~3�������uI���]� U��V�^�F9\sKK�9\v�\^��]�U��VW�N���w�F�( s!��r� s3�9�t�v�����uЙ_^]� A���S��w�_
3��#��[�uBS�w�_;�t6K3����T�;�s��r#��t���H;�s#�r�Э�t�����D����[�G�G��[�L�t	�+�H�+����ƌ���U�]�U���������������������� �>�������6��>� t� ���� �>�t&�>�t�>�t� ��� �>�(|h2 �e��E�F�t�>�tP�Nh �c�~ t3�P��� �� h ����:�t
��2��D����3���:�t@P�	��:�t��!���� ���>����6�� ��ø ���<u"��tErO��v������wK���D��+��������� 
�u+���$�$0<0t������� �� �� �������>�<u�� �� ����� ��� ����� �@ ��&�J �����>�|�0*��9���� �>��+����U��>�}� �F�>�|
<~<+~"�@����>�tN��0���� �����<��*��>�t.��0���� �������1�>�uԸ�0��� ���*۴���� ���>�th ��� ��C +��� U���<|/<|�2��^�e�����@ ���e &��~ u$�� &���� U����3��F��F����F������F��F�P��&�� P����t0;&u;$���;$~PQR�ZYX�#�&����������U��F�V� �����F�&�&��># t�B�� U��V�F�V
�N��r#���&��v�&�F��Iu��># t�	^��
 U��W�F
�V�N�U�r���F�&�����># t��_�� 3����U��F���� U��F�t������  �� ������� U����~ u�����>� t�������� U��V�F�� �>������ �$��;|%��;G�&��;G|��;G
S�?[�#�����r-�G��O�_��+��&������+ʋ�3Ҋ���ߎ����U��VWU�FP�^��X�N��tڋ͋���># t��]_^�� U��VWU�^3��fP��X�&�I��u�N�tڋ͋���># t�]_^�� U��^�G+G�W+�������� U��VW�^���W�G+Ћ?�&�������O+ϋ^��O�WU�������ێ�2�������J��tË͋������]�># t�_^�� U��VW�U�^����?��O���W2�������J��t������]�_^�� ��O+ʋ�W+W+��&�����3��������U����VW�^�0��F����~��F��G�&��������v��ߋ����J�^�����v����t�����&�� �V����J��t^�����># t�!_^�� U����VW�^���F�N��~��F��G�H�&��������~��ߋ����J�+^����+v����t�����&�� �V����J��t+^�����># t�_^�� ��>�� ���          ���&��t���5�!�������%�!�/5�!���t�D�5�!.�.����%�!�	5�!�����-�	%�!� ��r+
�u'&�Gt �5�!.�.���%�!� � ����%�!.��%�!���	%�!�>  t.��%�!�Ϝ.�.�.�π�OuPSQR����2��ZY[X�.�.P���؀>  u�`2�SQR�� ZY[X���.�> ug.�PSQR�&�.�t6�&�Ĝ.��&�.�t�&�̜.�� �Y V�о �  ^뾀> t
� �� ZY[X.�ϡ������؁��I@��;�t�  �w�W�O�G  ���<�t!��t�8'tC�? u�
�t2��
�u����Ĵ�P�&�Ĝ.�3�$�Ȁ>u��
t��X�<8t	<�t
�u�V�� ���V�� 3��Z�^� �35�!���t3��3�t�  ����� � �3� �3��"À>" t
�! �3�" À>" t
� �3�# À>" t� �3�U��>" t�V�N� �&�$�����3�� ���۩ t�  �=� t�  �(  �*� t�  �� t�  �� u�� �  � �����$�&�>+ t�> t�� �+ �� �> u
�>* u� �&�3۩ t��� t��� t��� t��3�PjSRQP�6 SRQ�> ut�&�&�_����;�rGw;�vA�� ;�r6w;�r0��6�;u46�G;u*��6�G ��{�(  �{�+���6��6�G��{��
��  �غB�$%�!�S�����Āt�݋\�ǀ�	u��2����[ϸf�!��s���U��	D�^�!r3��� u@�� ]� 3��2�t������2�ø@ ���&�2�À>D t���/�U�� �>D t���v�V�/]� U����W�^��^��G:\�G �ӌ؎��~� ��q��!� s3��,����_��]� U��V�F�v�u� �!����@��D:\��� G�>, t�Gq�!r3�����^]� U��;q�>, u� ;�V�!r3�����]� U��V�>, t�lq�^3ɺ �v��=�F�V�!r�^�3�^]� U��V�>, t�lq� 3ɺ �v��<3ɋV�!r�^�3�^]� U�� Z3ɋV�!r�^�3�]� U�� >�^�!r3�]� U��V�V� A�>, t�Aq3��!r3�^]� U��W�؎��V�~� V�>, t�Vq�!r3�_]� U��?�U��@�^�N�V�!r�^�3�]�
 U��V� C�>, t�Cq� �!� s3�����]� U��VW�~�>, u��>P�v�v�� ���u%� ��N�V�؎�� �Nq�!r��i3�_^]� ǅi��_^]� U��VW�~��i�u��>P� ���u�H ���i�؎�� �Oq�!r3�_^]� U��N�.�G��^��i���t
���t��q�!����]� ǅi��3��E��S���X�E ��Z�E"��\P�E,P����U��O�V�U��N�V�/�!��!<Nu�V�N���!P�P�ڋӴ�!X�Xr3�]�U��V�v�
�t��
u���!���!F��^]� U��F�
 �^�3����0�C�u��΋vK���D��D;�r��]� U��^� H�!s3�]� U��׋��v�~3�������+��t�������]� U��׋��v�~
�N�/��;Fu;�v���;�s��NO������ t�I�������]�
 �t�������� ���3��U��V�^� ^� s3�]� U��V�F�� ��^]� W�Ӹ =�!r�؉�� �� >���!�r_�_��� � ?�N�!r@�N=MZu8�T����f��?v��� ����3ɋ��3ɺ@ ��
� r�T ����QR� B�!� �?�N�!r;�u�Y=NStZY��&ZYS�P��� (+�[x�N���؎����?�!r��������3�&�ǉ������WU� ��]_�VS�( �h��<��� [^Ã�&���'t;�t����&}2�&�G��3��� U����^;�r� 	�1�> tO�F �tH�~
 t3ɋѸB�!rK�F
 uFVy(� ��6�V��F��ѸB�!FVy�N��V�� B�!�؋V�N�F
�B�!r������ U��׋ތ؎��v�~3�������+��t�������]� U��֋v�^��
�t,��'C8�t�,A<ɀ� �A��,A<ɀ� �A8�t������]�����U��VW�v�N�tB�G�t��FQ�I Yr	�ƀd��Y�8SQ�+�Y[Y����t���؎��WV������YX�� 3��Q��Y�V���Y3�_^]� U���VW��F�  At����INN���P$����;�sh�rZ��t�B�H����uA�Gt;�E�s�F� +��;s�RV�2�^Zs�F� ��r��� ����u��른 NN�#Z��9FF���F���t��u�FF�r�+�J�JY����%�	�W;�s;�v���_^��]��  V�v�v�j �F��uO�F�Pjj�dt�t-�F�P諤�u"�� ���DWh��6�F�P��u�u�^���t�A�>� t���7�j�v��tV藲V�7�[^�� ��  WV�^�7���uh��h� ��[�^�7���v�v��>�Pj ��F��^�7h�L�K���>�L u
j h�L���h�L�c��� �>� ��%2 Pj�6�6��6��oi���t� �>�*r	h�	hJ�&�=6���t� �^�7� �_���t� j ��6�K��I  ��>��"�4�t�t�#���tW諱��Ht��u��k~���>�;�w҃>B  uj j j j �����t	V�v�� �"j j �DW���B �r�6DW�2mj�1u3���Xg�;6�Zi��^_�� � V����Ph�Lh�h��_����P�g��tp����Pj �F�P�F�P覭�uZ����P�v�h�@h� �N�Q踮������P�v�藮�u3�~�� u,�>�@A<u$�>�@�Ru�>�@v�6�@��@ ��@� ��@�E��  ��@A<��@�R��@ ��@  ��@ �' �APh�hA�n��j'h�hTA�`���> t�A��TA������Ph�Lh�h��^����P���t����P�(fj h�P����Q h@h�R���^�� = s� ËЃ�<v�< �� V�>�  u3�^�Í���Ph�Lh�h�^����P�F�P������u����P�v�h�@h� �ح������P�v��_���^���  WV�v� � ���^��?/t'�?-t"kFF;�w� ��� �D�� �D��� �0|.�9(�GP��[�� �u�&� ��a=�v�� ��� �O�G�P�<�[=W t<w,Bt,t,
t��t"�G j ��[�$� ���  ��� ��,  ��&� �G9~
~�?���+F� ���^_��  WV�,�V�U�hD�O�GW�Z����< u�^_��R  WV�~��3��8k���F
Hu� HHu�Hu� - u�Hu�Hu��- u��Hu��Hu�- u�- u��-> u� Hu�'-M u�,Hu�2Hu�2Hu�2- s��- w�(-<u�)Hu�����3���j�V�߸ �j�M��v��u�t5�F�PVjB�N��^��*�Gk���"Kthw�`�P�F�P�n���F��EWjj j j �s�u�}t2�E*�����@P���6��u�u
j���j�6��u�EHPj���j3���.�v��>� t��v��Ru�FtW�v�jj ��F��1�t	W�v�j.V��� r��� wW�v�j���F�  ��Rt���~� t�v����WV� j���E�u��e�߸ �oi�� W謝W肞�~ tj j �֋^����m�E W�3lWj ��kWV�~	�[j �8��SWVj ��)��F�  �>� un�]�F�V��p�t)���bpWV�v�v�9WVj ���Ƌߺ �XWV���E��E9Ft�:�= u�
Hu���#pWVj(j ���F��u��P�����v��E9FsWVj��E9FrWVj��F9Ev	WVjj��9Ev���WVj��9>�t�3��oWV*�DDP�D*�DPj�x�g9>�u�]�F�V�p�u�NWV�v�v�_�D*�D;Du��D*�D;D
u�WV��!�v��>� t��v��u�Ft	W�v�j����1rW�D�P�<���W�v�V�v����v��vV��� �v��vV�7�� WVjj �� � WVj��WVj��WVj��WVj�v�ߋ߸ �wgk�v���֋�3��}g�ߍF��uf�F�*F��D�F�*F��D9>�uWV�Xj�?�j �w�߸ ���kWV���!�u/�vj�v�v�v�p���M�W�u�E W��iWj �i�!��vVj �D*�P�����v�v
�v�v�v�Fp^_��
 �  WV�~�v����ƴ �G*�k��� K�N�k���"Kt�Dt�# ���^�>�  t�Du� ���Dt	�v
Wj �T�v
�v�v��^����F��O*�k�9� Kt	�v
�v���Dt�v
�vj �y(��^_��  � WV�~��Fu4�^���u�؉�]�G�]�G$�>�I���= ��]@�G�3��t�*�Hu�]�  �]�G �]�G ��]� �]�G  �]�G  �6B �F�  ��t��YP��[��;~�v�F��4�u�v��6~��[��OO�6����[HH�F�ƉF�;�sI����2r�1 ��+v��v�j2j ����Q���߃�+�Ƃ�� �F�  �v���wk�zP����P�i F���뵋6B � �I�t�?Y�F�j2j ����P�j߃��v��s�[P�v�����P�(߃��^������� k���zQP� �4G�u��^�^_�� �  WV�~j4��[���E�F���D�E�vh��v�P����^_��  U��WV�~��u'3�k�zP�" F��v� 9uvk�zP�
 F��^_��  U��WV�~�uNN��EV��[^_��  �[��d
�u�& � j �l3�� j h^j h_j j �ǒ3�� j� 3�� ��  WV�V���u� R�9]���=��u� P�I]��
�=��t}�6������
�r����
��E*���1�w�����ލO��M�>1�u!�y��؋Ƌ��E��G����F�P�$]�F��%�'�h���j P�}o�������\���uj hhj hij j����^_�� U��V�F
=� tmv� ,t,�t2�w�N��-Grm- v
- rc- w^Q�v�v�^3�� �v3���Y���7�v�t�GP�\�D=��u�D  �� �D
�\�͋^���wj j �^3��� �:v�v�v
�v�v�v�o^��
  �  WV�v�^�w�h����E�D�E�^���G����u�H�؊�G�D�G�����<�u�^_�� �  WV�F� ��*�F��F�P������u� �6�����DW舔�t�B�!j j j��h��<����t�V���DW贖3�^_��U��WV�v�^
�F*G�D�F*G�D�*�Gk��� K�DD;�w
��*D�ȈD^_��  U��WV�~�} t!�v�*�Gk��D�� KP�]�T�� ��e^_��  �
  V�v�*�G�F��L*�L�N��L*�L�N�k���"Kt&�F� P�v�Q�F�P�F�P�?�u	�v���� �3������v��v�V� ^�� �T  �~�t�>F � t�F�� ��F �F��v�F@P�F@Pj �v��F�P�.����F�h�P�a���  U��V�6B �V��t�4J�u��tj j �֋^���e3�^�� �  WV�v�  ��*�D�D�>DW u	3��F� �� �F�  j h�+Vj j j jh�j W�'\�߉�DW�u����E�~��V���ڃ�DW t1�|u+�D��ڋ�DW9GwH�F���*�F������DW�F�P� �F�^_��  U��V�v�| u�LV�]�| tV�v� ��tj � b^��  U��WV�~�u�e��tV�^^_��  � �j_= ���ۋ�DW�V������u3�^Ë�3��G_^� U���v�����  �  V�v�  ��*�DjV�F
 P�gك�jV�F P���Uً^���G��O3���^�F��^�G*G�^��G8Gr�^��G�ȈG�v�v����j�v�.��v�a�vj �:a�^�G�uS�v����^��  �  V�v�-��F�=��u� �:k��^7���D  �D�D2��D�D�D  j j ��^�۸���DW��b3�^��  �>DW t�>FW t� ø ��  ���Hu&�F� ��*�- �+���@@�F��v�v�F�P�d��3��� �
  WV��= uJ�^����]���F� ��*�F���������DW�F�P�^�����3���DW���^���DW��\W�)\�D3�^_�� U��V�v�������tV�\3�^��  �t  WV�F�  �(�Hu�>� u3����F�  �v�F�� �*�DW�u�É^��6FW��FW�F���>��� �F��|�~��F�P��j �v��Ր�v��_j ���v�VWW��v��~����~��NwL,t	,u� �?�F�- u� - u� --t- t
���vN���*�- ;�vFW�v��v�V�>�v��F�P�Ta�F�= u��F�+ҋ���s� ���*�;�s���t$��wj h� ���*�;�wj h� �j h� ��9v�t�똋v��~��3��c��w
Wj j �1��z��*�;�w�u�F� �T�v��ރ�s� ���*�- ;�s
��*�����F� �v��u�v�v�F�P�9��F��#�v�W�F�P���F��F��*�F��v��F�P�s���  �� ۃ�DW u�>� ��أ� �� ���DW�Z�� ���DWj �4^�F�P苏�F�^_�� �  WV�^�v�G*�����AP�7܃�v&��*�;�v�6�Vj j���[�6�V��*�HPj���[�v��vW��*�;�vN�6�VjjĠ�HHP�0\�6�Vj j��[�6�V��*�HPj��[�6�Vjj�[�6�V��*�- Pj�[�~
 u1�F� �F� ��*�H�F��v���v3�6��F�Pj �^�GP��[��~
�u9usW��3��lZPj �D�P� �D�^�G9Gv�^S3��KZPj ��*�+�HP��^_�� �p WV�vV����P�у�V�N�u����P�v�6� j �����N�~����PWj�֛���u2����P����Q�EM����P�v�vj ����u����PW�ޛ�t�3�����P���^_�� V�6B �tV� �u�4��3�^ø ^��  WV�~3��E*�k���"KtVj��4���uK�uj h�h�B�睃�j h�h�h�Bjj��"��F�Hu� ��~�uj �EPj!j �d���tV�|���^_�� �  Vj j j �F�P�� ���uj j �^���V��]��^��  �  WV�~3���F�P�D��t� �>D uPPPP� ���tV�=a�t�vWjj ���^�F����t�9F�u�^��PVjj ���B 9F�u�^���B ����؋~���9?u����E*�P�!���u��[W��[�>D v�D ��^_��  � WV���F��>D 	u�" �]�~
�uG3�FVj h|����P菜������P�t�u�N�F�  �~ t,����P�Y���t�^3��?�����PW�F�P�,J�u��� j-�7�[�F��u� �� ����P�0�[@P��[���u	�v����[�܍���PV��΃�j �V�~
 u:�v��F�=��u�F� �~� t� �D �^��w�F��G�  �B �V����V����t�V�F�P�v�v��*�F�뾋4�< u��~�F��؉�G���G  �G�G�G �G�G�G  jS�GP�5у��t�F����v��/�[V�*�[�v���U�F�^_�� �  WV�v���F�j ��U�*�Gk���"Kt�vVj"�v������w�G*�P��-���u�*�Gk���"K��v��U��^_�� � WV�v������S3��F���S��S��Gk���"K��S�t��Q �#��wh�P�t̓�h�P�QJ��Ph�Q�b̓�� h�V脘j ����P�.�h.j h�P�b�t�� �tHu�� @@u�� � �������G�*�Gk���"K��vVR����F��t���S�O*�k���"K�v����F� �bW���[����PP��[@P���[��P��̃�j W�^� ���Y�^����F��t��^�9uj W�^����ظ ���Y�*�Gk���"K����~� t�"��~��	�& ��>B����P�|H��^_�� �
 WV3�h�V�p�V����P�ލ�����S��S �6�S�~h�	j h�P��`�u?�t	Ht>@@t?�2����P�6� �6� �F�P�a����uj j �߸��V�� Y�V�ؗ� �u��	�& ��6B����P��G��^_�� �
 WV�~��3��JT�F��F
=� u��v��,t',mtJ,tc��u���u�,0u��,u��W�^��� t�j ��� P�v�v��h�t3����^��� t�~t�kW�v�9�a�~ux�v��^������؊߁�� ���W��ȉN��V�RQ�*  ��������P�v��v�W��ƃ�� h� ����j P�^� � �gj j j �^� �� ��f���v�hr�I��F��vj j �^� �� ��f�؉F��[uhF�v��Ĩ��^����A*�Ph�hH�@Ph�hL����P�{����� t����PP�� t�����Wh��Dh� ����j P�^� � �cfj j j �^� �Q�j j �߸ � �3W�+�^�v������Ë���ˊ߁�� ����x���^щW
�WR�*  �^���G�b��v�֋�3��YRh� �� t������F�j P�߸ � ��e�� tX�� % Pj j �߸ �� �e�� % Pj j �߸ �� �e����P�6� ���h� ����j P�߸
 � �xeW�� % P�+V�;E�t����j V��ڍ���PV��Qh�CW��V�aWVjj����P��W�v��* �u���F�P�YI�v�v
�v�v�v�^^_��
  �
 WVj j j �^� � ��d���< uj jPj h�j j���������PV�F�P�yC���u��Ht- s��- w�� ��v�� u��t������P�߃��uj#�����P���ȃ�����P��D��P��P�ȃ�� ����PV��ǃ��� ts�&� �j j j �^� � �%d�t�� j j j �^� � �
d�t�� j j j �^�
 � ��cP�I�[�� = s��  � �� =�v��� ��������t�j jPj h�jj���~Hu��� �~��v�׃�u����PP��Ph��A����P���,ǃ�����P�D��� ����P�8C�F��us�~����CP��P��ƃ�h� ������ t������F�j P�߸ � � cj j h������ �n �c����Vjj���V ����������P� �v�蒒3�^_�� U��WV�~�v�޸ �c��W�v�D+D@P��j W�޸ �� �S^_�� �  WV�^�F��b���^�F��b�F�W�v�F
P�D���v��v��F�u���tV���EuW�QWj�.Q�v�j�&Q��^_��
 U��WV�^�v�	 ���gb�؋��>N�߸
 �Xb�؋��/N^_��  �  WV�~�v�F�  �E�F��*�Ok��� K�;�s��+F���ƉF�+��v�~����~� u�v
�vW�F��P�9 �F�GN�u�v��v�N����v
Wj j �^*�GP�OGN�u�F�^_�� �`  WV�v*�D�F���GP�v�F�P�t�v��/=��u� ��| u�� �^����DF;F�r�DF;F�v� �|�F�;�sL�v
*��\��P�O�V�vj �F�P�F�+�P�:N�F��;F�v=�\*���GP�!�9~�v�F�+���v
��3��F�V�vP�N��P�F�+F�@P��M�F��;F�v`�\*��Ƌ6��Q����͋F�@�v�;�v�F�+�@�3��F�V�v��P�B�PjP�"�^
�_*��6�� P���v
�vj �F�P�v��M3�^_��  V���| u3�^ËL9Ls�L�O�L��O�L�O�L9Lt�O�  �G � ^ËL9L
s�L
��LI�O�	��D
H�G� ^��
  W�^��F��Hu;�V�F�+F�@�F�;�rJ�V��^�*�GP�v��v��F�P�v�*�^��~� ��% _�� �  WV�v�F�  �^
�G�F���ÊV���^��^
*�GG;�t/9wv�w�*�GGH;�s�ƊO*�+�@�G�^
��*G�G�^
�V�G*�G;�tH�G�F;�v9�Fw��+�F�#3��*�GG+�FH;�s*�G+�F���@�G�^
*W�W�F% �^
����F�u|�t�v�v
j �^
� �F��^
9Gt� 9tW3��F��F�G�F��G�F��v*��\�6�� P�ˋ^
�G+�Hu+�v�F�Pj�fL�v�^
S*�G��HPOIQ���:�v��7�G+�=��u�v�F�Pj�SL�v�v
j �^
�w���vSj *�GP������^
9t�^� tj j �~
�_�U�� �N�v�v
�/��^_��
  U��WV�~�׃��^�F���d �^�F�G�F�G�F
�G�F�G���~ �v�vj �^*�GP�`����^� tj j �~�_�U�� �BN�v�v� ��^_��  V���| t��u)SPj �g ^���t�D �D*�D�D�D*�D�D
^� V��| t4�t0�D*�D�D�D*�D�D�D9Du�D9D
u�D  � ^�3�^� U��V�v�| t�D  �V�tRVj �D*�P��3�^��  U��V�v�v�D*�P�DP��JV��^�� �  V�v�D�F��L*�N��L���Ok�9� Kv�~� t�N��F��vV�t�D*�P�v��v��v�l�^��  �  V�v�D�F��L*�N��t�D��*�;�v�F��N��vV�t�D*�P�v��v��v�"�^��  U���v�^S�w�G*�P�v�GPj �����  U��^*�GG�@�O*�k�;� Ks"�v�^S*�GGP�G*�G@P�v����3���  U��^*�GGt�vS*�GGP�G*�GHP�v����3���  �  WV�v�*�Gk��� K�D�F��L*�N��L�9� Kw��*F���*�F���D*�F�F�;�r
�D*�+��~��vV�t�D*�P�v��v��v�
�^_�� �  V�v�D�F��L*�N��u�F���D*�;F�r�F�  ��D*�)F��vV�t�D*�P�v��v��v��^�� �  V�v�D�F��L*�N��u�F����*�HH;F�r�F�  ���*�HH��F��vV�v��v��t�D*�P�v�W�^�� �  V�v�D�F��L*�N����- =�r��*�- �F��$��*��HHF�N�II���v��*�- �؉F��vV�v��v��t�D*�P�v���^�� U��V�v�vVj �*�Gk��� KHP�v���^�� U���v�vj j �v�����  U��^���u�B j j �ы^���+J3���  U��WV�6B �~�tW�t�Sԃ��t�4����3�^_�� WV��= vG�� �3���DW�?E���>� u3��� �3���DW�$E���9u�D�� �D*�DH�� ^_��� ����   ^_��  WV�V��*�GG��;� w-9� w'�>� ���ۋ�DW�^�3���D���v�P��+EPV���^_�� �  �>� �tt�� 9Fwl�>� ���ۋ�DW�^�3��D�F��� 9Fs$�^��V�G*�G� �+�;�sW� � ��v��v�j �^�*�GP����^�� t	�v�Sj ����  �  WV�>� �t�� 9Fv� �~�>� ���ۋ�DW�^�3���C���F�;� s)|�/�*�Gk��� K�F��L*�L;�w9|s��D  �F��ȈD�D�� �D*�DH�� �D  �v�Vj �D*�P�+�^_��  U��^*�GG=�s�vS*�GG@P�G*�GP�v���3��� U��^*�GGt�vS*�GGHP�G*�GP�v�Q��3���  �  WV�v�| t�vVjj �8܋��us�D*��|�DD�F��>< u�*�GPW�v�j� �F��uA�F�F��*�GPW�v��F�Pj�^�u!V���vV�F�@PWj ����vV*�DPW��^_��  �  WV�v*�D���|�GPW�DDP�F�P�!�F��u)W�EPj�����vV�v�Wh ��e��vVj �D*�P���F�^_��  �P  WV�~�F�  �*�G�F��M*�M�N�k���"Ku�^���]�= t� �6�@�B� �FtQ�v��~�9v�rl�~� uf��@�F�WVj �F�P�F�P�] �F��u!h��F�P�&���;�@rWVj �6�@�l�F�F뵋v��~�9v�r�FuWVj �F�P� �F��uF���v�vj �^*�GP����v��v�j ���S�FuM�vVWj ���v��E*�E�F�P�v��F�P�4 �F��u#W��VW�F�F�P�v�j �$�VW*�EP�v���F�^_��  �  k^
��"Kt�F�	�^� �F��F��V���F+��6�@@�&�@�^+F�+��F��F��v
�v�v�v��v��^�7�6�� U���v�vj �^*�GGP�v����  �  V�^�7*�DP�GGP�F�P� �F��u�v�v�v��^*�GGP�v�L�F�^�� �  WV�~�F�  �*�G�F��Ǎ^��j��tHu� Hu�� �!�E*�E�F��E*�E�F��v��v��F�P��F��t�� �F�9F�rBk^��� KH;F�v4�v��v��v��F�@P�u �F��t�� �vWP�E*�P��F�P@Pj� �v��v��v�j�B�F��vW*�EP�v��y�W�M�W�����v��E*�EP�v�F�+F�@P��F��vW�v�E*�EPj �=�W���G�v��~��W�v��|�F��u1F9v�s�v��~�vW*�EEP�v�j � ��v��v��F�+F�P���F�^_��  �  WV�~�F�  �*�G�F��EE�F��M*�M�N��t>�v�Q�F�P�]���t� �vWjj �׋��u�F�9F�v�~�vWjj �׋��o���t�v��D�P�F�P��F��t�T�v��M�v��F�HP�v��v������u6�~��v�v�v��E�Ph ��F��&��v�vj �^*�GP���v�Wj����^_��  U��� �F � �v�w�3���  U��� �F x �v�[�3���  �  WV�v�*�G�F��DD�F��D*��|�v��v��F�P�G�F��u/9~�v*�v��v�W�F�+�P�G�F��u�v��v�W+~���W��F��vV*�DP�v��O�V�#�V��ۋF�^_�� �  V�^�7*�D�F��G��w�v�VV�P�F��u.�v�V�b�F��u �v�vP�^*�GP�b�VVj���v�qۋF�^��  �, WV�~�*�G���EE@�F��F% = �@�F��F�Ph���"Ɔ�� k��� K�F�E*�E�F��v���v�9~�w�� �v�W����Pj h��4�F�=��u� �~������V�����f�~������*��F�؀��� ��"�*�= �@= ���;�u5�����;�r)�����*��F�؀��� ��"�*�= �@;�tF��F������;�s��~�G3��S�� ��v��v�v�ƍ���+�P�v��v���3�^_�� �& WV�v�*�G�F��F�Ph���!Ɔ�� �D*�D�F����{9~�u�^*�OO��ȋэ���ЉV��~����H���*��F��*����� ���u)����;�r!���*��F��*����� ���u1N��N����;�s��t>O�v�W����Pj h�������t�j�� ��v��v�v�ƍ���+�P�v��v����3�^_��  �  V�v�^������HtHt �% �,�*�GP�v��v��F�+F�@P�X��*�GP�v��v��^�� �  WV3�96�Iu3��� �~9ut�vWjV�WӋ��t� �>�IuP�K3�����V��u� � �*�GP�EEP�E*�EP�N��DQP��&�4��F��K3���W����K�v�kK�� KH�F�3��~�!�*�GP�EE�P�6KV�E�F��uF9v�wڊE*�EPPV����vWj �E*�P��W�؋F�^_�� U��V�v�vjj �ҋ��u�v�vjj �lҋ���^��  �>K�t�6K�`3���IP�c�K=��u� �3���  Vh��x�[�F��u� �I�����u7�v
�v�v�FP�v�����u�6Kj �v��vj �����u��I �v���[��^�� �  WV�k��F��u+3��v��6KW�vV�1�F��uFG9vs��t��I �F�^_�� �  WV3����F�Pj��f����~��w� �x����P謴[��S�u� �h�~��v��6�S���tV芴[���t߉~��>@W�BW��D��P�?ċ��u� �*�@W  �6BW�v�������u�K���������Kr�3�^_��蕡��  WV�K��<�t	�����Kr���Ktj ���������u� �������S�G���@W�&�G  �@W�&�G&�j 躡�F�=��t~�����S��������S���S�����@W�&�G  �@W�&�O&��F� �F�  �N�QjjP�� �t�v��Ρ� �D �F�D��-K� ���P���r ���	W訡����^_��  U��WV�~9>xu�z��9>|uj ��k���K��6�S���+�S��P�`�����S���<�u�k�ǇK��3�^_��  U��V�^k���K��K���6�S��؉O3ɉO�O
�O^�� �  WVj苠�F�=��u� � ����F��V��u�v�����^�Ë^����6�S� �����Ë�S�֋H���H�����>�S�N��	��S���I���>@W�N&�	�@W��� +F&�A�FF
t�v��v��v�v
�v�F��ן3�^_��
  U��WV�V����6�S9zu��z��\���>�S��D�4��S���@R�!�^_��  �  WV�~�����F��V��u� �W�����@W� &+I��V�ً��~�&���^&�]�]S�v
�vR�����r��@W&��@W�F &)A����3�^_��
 �  WV����9Ds+D�\�( �9|v�D�\+��� �F��u�|�F��3�^_�� �  PSWV�O��G�F�N���N�����@W�BW&��F����;�w*�����6�S�����8�t��+F�ȋ�3��~���� �[�N��~�������F��V��u� �A�v��^�N��~��G�v�&�  �I�u�~��^�F��~���%��u�F��E�F�E3�^_���  PSWV�W�O��;�s9����>�S�]�}��>�S�}�t��@+��^����>@W&�	I�V��ȸ �h�V��v�N����P��F��V����u� �I�~�F�)F��F��F����F�&� ��N�~� u�^��F��~���o��u�F��E�F�+F�E3�^_�� �  WVk���K�ߋ��2��t3����E�Μ���V��t�EƋV�^_���  k���K�^�������u	�^��G������  WV�F�V�����V��u����>�N�F�&�5;�r��N�v
�v�EPV� ��~ t�F�&�E�^*��F�V����^_��  �  WV�>�  t��>�  t� �Lj�{���uA�F�V�����V��u� �*�v
�v�N��DQP��&�4&�D*�P����F�V����^_�� U��WVk~��K�>� uj����u6�ߋF������u(�v�vj �F ���u�v�v�v
�v�v�v�����^_��  U��Vj�����u�v�vj� ^��  �  WVk~��K�EH;Fw�.�~��ߋF�y����t����~��E�F����F�V��u� �� �v���6@W�BW&���uO�~ t)�]� �m����t��u��]� �����u��v��O��^����6@W&�   ���@W��&�@ � �E�F��G�;E
w,�]� �����t��u�]� ������t	�F��ƚ�@��^�v�&�  �F��^����>@W&�	���@W���N�&I�V�^��SR�SR�@W�� &+H+N�Q趼�F��p��^��O�O3�^_�� U��V�vVh���DPh0��< t� �3�^��  �  WVk~��K�} �r�$ ��~��>� uj����t���� �^��F������u�v��~��E�F��M�N�����@W&�@�F�N��;�sW�v
�v�v�v� �F�� �F��C��V��u� � ���v���N��~�N�~�EQPQ�v�� ��+v�V費�F�^�&��N&�O�OQ�v
�vP蓻�^����6@W&� �F ���@W��&)@�F��.��^��G�~� u�^��O�F�^_�� �
  WV�F� �^��w��蔘�F��V��u�� �v�PV�^�w
W�_��F��t�� �v��F� = vj j j j W�9��F��u5����S���@�F�P�v
�v�v�v���F��t ������S�p��������S�p���h�v�ߋD
�����>@W&)�F����@W&A�v��^�S�V��RS�@W� &+QR���j����%��F��D�F�F = v3��D�D
�D3��������F�^_��
 �  WV�>z�u)�x�>xr�x  kx��K�t�kx��K�z�z�����S�7���u�� � ����@W�BW&+G�F�� ����@W&+O�N�&;Gw�����F��V��u� ������F�V��tpkx��K�^�9wu�F�G����@W�BW&��^�G
��F��V�F�RP�v��v��v��O����@W�F�&)A�������>@W&�	��&	V���6z�z����6z^_���x  �z������>x u��>z�u��U��WV�v�~���ЈG�< u�^_�� ��  WV3��F�F�F��F�  j����t��F�Ph h h���F��u� ���v
�F% = �% P�F�P�F�P��k�F��t��9F�u�Njj j �v������
������u� �v��� v�F� �vj j j �v��չ��j ���=��u�F�" �ek�K�؋�����S�������@W�BW&�  ����@W�BW&�G �E  ��:�P�@_j �v
j jy�F�P�o��
�F�h�P��^�F% = ��؉F��t
�~��F���~��F��B�F��F��~��F���9v�ul�v
�v��v��v�F�P��k���t�� �v���F�F��F���
F�kF�
+��v�k�
�F�;F�v'=d v�d �F�P�v
j jy�F�P�o��
�F�h�P�D^�<	u�~� t��+��6�@@�&�@���G�~� t9~r�~� t�<
t��^��F���d�F�  �~� u�~��Bty�~� t%9v�v�<
uF��F� �~��Bv�^���u�N��F�-�BP�v��� ���u-�^��G���s%�F��B3��~� t�����v�^�7��� �~���j(�m�Nj j � �F��t�^�7���~��E�^�7�1�~� tV�}vP�^��F��UJJ�V��j����V��t4�F�&�<u&�|u�F� ��F�  �F��V��t��~� t	�v��v����F�E��:�P�G]�v
�v��*j�v��t�[�F�^_�� U��WV�~�6����@W�E&9@s:j j j j �����S�7����u+�>�  t� ������6�S� ���6�h�BW�v�m�^_��  ��  WV�~3��F�F��F�  W�'��uW��u� �pj�����t�`�F�Ph h hh�X�F��u� �Eh�¤[�F��u�+�vP荟�^����G S�F�P��h�F��t��k^��K��K���6�S�0�N��؉N��O������ىN��F�  �O�N���Ñ�F��V��F�u� ��v�8�P�[j �vj jz�F�P�2l��
�F�h�P�e[�~�v��F�H;F�w��F�����BW@W&9w;�F�  ��輑�����S�?�����S�?�u�� ���6��F��V��F�u�� �^�&��F�@@�N�+�N�;�sp�v��v��v���+F�P�h�F��t� �v��F�
 +���F��u�F� �F�+��v�k�
�F�;F�v'=d v�d �F�P�vj jz�F�P�Ik��
�F�h�P�|ZV�F��V� RP�v��1�v��~� t�^�&�Gu�F�
F�F� F��F��F�����v��v���v�� �u�F�9F�v�v��v�P�F�+F�P��g����8�P�`Z��艐�v��v��>g�t�v��nh��~W�eh�v�W�th���v��l�[�v��e�[��^_�� �  WV�V3��tR�j�[�F��t%�v
�P�Y�[���u�F)�9Fv��v���[��^_�� �  V�v
96|u�HW9Fu�^�>W��^��B�_�,�ƋV��V��u� ��؎F��v&���v����D3�^��  U��N9|u�HW9Ft���V�p��� j � �U��SPWV���|9F�u9HWtQ=��tj�e ���u[hj h�B�~����v�Wh�Bh h8W�B�>W=��u� �/�F��|�>HW3��~������9F�t�V����F�� ��3�^_��U��V3�96~t&9vt!���6|�6HWh�B�6>W�68W������|���~  ��^��  �  PW���B�F�k^���"Kt���$3ۿ�B9~�v�=	u��+��6�@@�&�@���CG���_��U��RW��k���"Kt��_��3ۿ�B��=	u��+��6�@@�&�@���CG9^�s��-�B_��V�6>Wj	h�B距���tCh �E�[���u� ^��6|�6HWVj h ��>WPVh�B���|���o���V��[3�^� U��k^�� K+FHu���v�vh�B�6>W�68W�~����3��� U��WV�F�V�^
�	����t����v�v�����u��@����u�F>W=�v�� �F�=�v�� �~�>W9�r� +�P���BP�F��BP�ۜ���vj ���BP�=����V>W���J�=�v4�>W+�P�F��BP���BP蘜���vj �>W�BP������P�>W9�v���>W�F>W�
�F��>W�FFt���BP�v�v�v�ˮ�~ k���"K3���I��  ^_��  �  WV�v���r	�-��  � �F
�V��������t��� �v
�v�a����u�������u�v
���B�F��VV��������B�+��PW�v�賛���~��>W�B;F�v�>W�B;�s	�>W�B�F��F�+F�>W�F�+F�Pj �>W�BP�曃��~ k���"K3�^_��  U��WV�~�v�v
�v�v�5�+�����u� ��3�^_��
  U��V�F�V3�������u�F�>W���^�3�^��  �  W�~�Nϋ�3���? t�?	t��C;�w��u3����+�@_�� �  WV�~
k���"K% �F��ǋV�^�i����t�Q���v
�vh�B�6>W�8W�F�P����t�(��;>Wv�>W�>W+F��~� t
�V��F�  �/�V���B��? t�?	uC���B;�w�^��Ӂ�B�F
���F��^�F���v������BQ�BP�����v�j h�B�m����~� uh�B�F�F�P����F��v
�F@Ph�B�v��v����F��u�v
�vh�Bh �F�P���=��u	� �R���N�~� uh�B�v�����F�@=�s�^�Ƈ�B�F��^�Ƈ�B
�G�F��v
�vh�B�v�j �y�j ��3��j ������^_��  U��V�v�D4 j jPh�Vj j���M^��  �  WVj�a����t� �F
�V�^����F��t� �~�v
�Ƌ����F��V��u� �|�N���&��F��=�v�Ƌ�����٢�  �Y*�&�G�8W���BP�GP�v��%��Ƌ����V���>W����=�vj �����~ VW���F��tj ���F�^_�� U��WV�v�uj���t	3��'�~�
�~��B� �v
�vV�5j �o�=��t׋�^_�� �  WV3��F�F��v�v
�F�P�F�P�5��t����� �~�vVj W�R���k^��"Kt5�F9F�v)F���F�  9v�v�v�W�F�V�FRP;v�v�v�V�%��q�F�V��F��V��~����~��J�FF;�vK�~� t�N��'�^��F�&��F�<	u��+��6�@@�&�@+�H�F��F� ��G;Fr�F��F�F�F�;F�w�+v�v��v�v
���F�^_��
 U��V�v�B  hlj V�4)�u�vV�c �B^��  �  V�^� u*�GG�G�G*�G�G�>�K u�v�v�v����vh�K�� ���u�v�v�	 ����^�� �  WV�v�D+D
��F�v��|v� �� ��F��F�v�^�S�w
�wh ��~Ћ^����G �vSj �^�*�GP���3���F��F��F��^_��  �  WV�v�|�D�F��D*�D�D�D*�D�DV�v� = t���� �|�F��D��^_�� �^ WV�v��~�G*�F�k��� K�F�} u� �Sj������t�E�F� �EP����P�咃����u����P��[������v�F�Ph�����(�P�ZO�D�F��D�F���9v�w� �^��*G��u$Vj j~��~�P�_����~�h�P��Nj�"�ub�v�Vj �F�P�����tZ�~� t�^�F�W����F���Ku�ߋF��-�^���F��P�F�+F�P�7�F�P�p �F��uF�F��f��& �v��~��F� ��~��v��v�D �F��D�D�V�+V��F�����D
�F@@P���[��׋F�����D3���(�P�yN��^_��  �  WV�v
�F�  �v�ȑ[�F��~��V
�F��;�vl�^���: uXG;~�u��FtQ;�v�L��������^����� ���t+�F��;�v#��������؋~����� ���uF3�닋��3�^_��
  �����?a|�?z�'�C;�w�� U��WV�~j j W� ����v��������؀����F�< u�^_��  �
  WV�~�E�F��E�F��E�F��E�F�h�j W�l%Hu�@@u�Wh�K�������&u��tV�f\�u͉v���Kt3��m�v�v�e��6J��؉F��G*��*��؋^,�O�^*�O;�v����*�����>�(v����Ƞ�*����*��^��GhFj j ��$�����u�� ��u�� �v��t� �^�?*�EP�w�w
�G+G
P�<����uoh?L�ڏ[���F��^�?*�EP�w�w
h?LV���F�=  u%h�K譏[�F��^�?*�EP�w�w
h?L�v�����u�^�G
F��G����v����u�vh�K������&t5��t0�t�v�v�1�V�[� ��Ku�v���t����6B�3��^�G  �vS�v��F�*�P�v��F�Pj �i̓�u� ���3���B^_�� �P  WV�~�F���fu.�t'�>@�u �6�  �F�P���u�F�P����6��^_�� Ȅ  WV�F
=� u� v�,t,�t��vhH �v�v��+�u�� 3���� �~h� �F��P��|�Ph� ���u��|����Kj V�߸ � �T*��K% Pj j �߸ �� �>*��K% Pj j �߸ �� �(*� �~j j j �߸ � �*���< u� �LVh�K謍��3���KPPP�߸ � ��)�t��Kj j j �߸ � ��)�t��K�6�h�K�������&u� ��^��W��tV�JY���v�v
�v�v�v�#^_��
  Ȅ  WV�F
=� u�� v�I,t,mt$,PtN�:�vhV �v�v�*�u�$3�3��/�~t��vj j �V��޸� ���K�ދF��V���(�� �vh� �v��|�Ph� �*��u��|����Kj W�޸ � ��(h� j h?L�޸ � ��(��K% Pj j �޸ �� �(��K% Pj j �޸ �� �(��vj j j �޸ � �(Ph�K�5���j j j �޸ � �s(Ph?L����3���KPPP�޸ � �V(�t��Kj j j �޸ � �<(�t��K�^+��G�� ����v�v
�v�v�v�!^_��
  U��F
-x u�~u
�^� ���'�v�v
�v�v�v�k!��
  �`  V���F���G�W�F��V���@���� RP�F�P�X���F���G�G��^��F�Uǋ��F�j ��B  h �F�j P���uJ�~� u�F�  �^�*�Gk��� KH�F��u9v�u!��@���� �^�*�GP�v��v��" �B�F���V��G�W�v���B^��  Ȱ  WVh��ˏ[�F��u� �� ��P�P�8Gj h� ��F�v
�F�P�S���t� �F� �v�~�9vrfj��uX�vVWPh����F�=��t?�����G
�v
�v�W�F�@@P�LT�F��uVPh� �F�P�GW���F�h�P�zFF럋v���& ��F��v
�v��F�Pj�T���v
�v��S��P�P�F�v��֎[��^_��  U��V�F
-� tHHt�8�v�^�?���FV�K&�6��vjj�m&����u3��� �^���v�v
�v�v�v�N^��
  �(  WV3�j'�6��F�P�G���hZ�F�VP�#�����u�6B�uj'�F�P�6������6�j�K��  ��^_��  �  WV�F
=� u�8v�,xt,t4,u�� �|�F- t�qj'�> t�����P�6�趋���@�~��HtHHtMHHtI�?�vV�F������F�P��j��F�$�j P�޸ �� ��$j��F����~j P�޸ �� �����M�F��> t	�^����^��*���6��6���u	�F�$����	���N���
��F�P�o�v�F�P�A� �v�~u
j h��t��> t���j h��\*�P�DP�~ �D
�\3���m�F���>�%  ��Pj j �^� �� ��#Wj j �^� �� ��#jj j �^� �� ��#j j j �^� �� �#�v�v
�v�v�v�8^_��
 U��WV�~
 u
�v�뜋���~�v�hPW����@�N�u�hPW����^�����^_�� U��SWV�����n�v��*�� ^_�� �  PV�> t������F�8F�u���+�^��U����F�G&j j j �^� � ��"��  �  WV�^ۊF��n���N��
��F��~�H�Dt�F���F�F��Dt�*��2F�$0F��Dt�*����2F�$2ȈN��*��F��FF�<'u�^_�� WV3��>�@h�VV��=��u�u�6B;>�@tj����6�j�)��^_� U��WV�F
-� tHHt0� �vh��6�@蓚h� j h��޸ � �"V��@ P�["�S�~j j j �߸ � ��!P�K�[��聡;�tj h�j h�j j���<3�3��,�6�@Wjj�F"- ��@� �� ���v�v
�v�v�v�.^_��
 �  V�v�o�[���t�v�v
�-��^
���@�<\t<:t� \F��+v��V�vF
P�T����^
�v�@� ^�� �p WV�~�v�vh������P�v� ��tHt$3�� �v�V�t� �s����% = �FF�c�v�ӄ[�^���@��F�<:tJ<\tFS��u��v�F�P�M��u��v�v��N����P�v�G �u�v����P�V �v�8O� �� �= u�v�vh�M��t�v����P�' ��^_��  U��V�v�vj�N���v����^�� U��V�vV�� ��� VV�vh��^�� �  W�~W��[�F��tV�e��F��}:u��P�Ʉ[-@ P�U�[�t.� �3�^��y�\u��v
�y�:t�A� W誕�t�v��%�[�ҋ^���u�3�_��  U��V�vhRV�0����؀8�@^�� �  WV�~W�F�P�cL���uW�v���L��W�N�����^_��  U��WV�~j\W踄�����uj:W�������u����D^_��  �  WV�~�v�~��v���FH�F�� �t�= u�� �}:u��% ���D:GG�3Ҁ=\u�u�7�@��D:FFG�~��~RV�a��t� V覂[��|�\uN�\�V��^�? u� �?.u3�.u-�\t� u!N�<\t�<:u��<:ty�F�^�? t��F뽀?.u"�\t� u�F�݀? t;�v�FF���^�?\u�;�vF�\�^�?\t�{��� �@�|�:u�\F� � �0�vj V蟓�t�FHP�v��v�������^��v�@� ����3�^_�� �r WV����P�vj��K���t��u�^�? tS��h�胆[�F��u� � �^���3����� ǅ �t� �~�v�����P� ���t]�v��~��>��� thv�j�����P�L����v�D�F��Lj j �޸� ��!j j ���޸� ��F��D�~�u�����PW�vK���t�뒉v�듋v��3�����P蝔��^_�� �  WV�v輀[@�F��^�� r�' � �� +�;F�sT�� @s�j�fs�� ۉ��� ۋ����tǋ���r�� ��� �P�� ���@ uW�s��� Ǆ  �� H��
���ۉ���� ���@��P��RP�v�v����F����3�^_�� U��WV�~�v+>���z����������Ê߀���� �>��	�Q�RQ��+߁�z��������Ê߁�� �	�Q���RQ�y�^_���  WV�^3��?���ދ��^��Cr�^�����rF9� w�W�<�[�^�  ^_�� �t WV�~�E�F��Mj j �߸� � �I�F��uz�v����P��~��h@����P���P��~������P����Pj�UI�F��ui�v����tH����.u���� t:����P��~[j P�����޸� �����t�~��~����P臒�F��E�~�uc�f����P�v�+I���t��~��~�e�3���sȀ��V t5�DA*�Pj hr����P�jK������P�e~[j P�����߸� �c�F��u�F뼋~��3���^_�� U���vh�jj �R��� ����� U��>��u����j �v� ��  �  U��WV�>��u����#�~�EPj�� �����u	k��� K��+�- ^_�� U���vj�v� �� U���v�F P�v� ��  �  V�F�x �>��u����%�6��FFP�v�F�P���t�^��v�  �F�^�� �~  WV�v�~�%�^��F��� P�= �F��t���t(P�}[;�tF�F�x �6�V�F�P�F�P�4��u¸�����^_��  U��V�vh�V��~����<@u�|@u�|!u�D�3�^�� U��>�s� u
�>�
s� �b��q�� �vj�U�j ��j j �a��L���>� u� ��F��t��������~
 t�`��tj j 贋��*䣂����@����h��j j � 7��P� �+�=�t��.3��� ��
  �?��>u�  �Z��l �Y��  �V蠂�>�t�>�t�>�uGh ��Ҁ[���tV覀[��*�@��*�����@ ��P�|����t+�PQ��RQ�6@袐^Ã>� t��+�PQ��RQ�6@腐��  WV�>> t*�v��HHt- t� ����?�V�u63ɉN��:��?��v�ދ�HF
" P�)�[�F��uj��F� ����ËڋO�G�F��u�F�E�F�E�F�E�E��^���M
G�E�GF��E�GF��E�Ft��t�E
@�E�EH�	�E
�E�E�E�E�E�E�E�Ft��t�E��t�M�~ u�ދ�^��F�E3��E�E;�u����~��ڃ���@@�؃? u��^���^���uj ���~�� tL�� t#�^��G�F��G
�F�G@�F��G@@�F��F���F�
 P��^��G �^��  uj��E� �J�F��؉G �v�v�^�� ������u,�Ǩu�^��*
�v���v�j��^��tS�' �F���^��  �>> u�v��b~[�6B3�^_��  �  V�v�T���Dt'�F�  �D+D�F��D+D�F�@�F�V�F�P��R� ^�� U��WV�vjhL��vV�DPj j �vj j ����j �u�ދи� ���^_�� �  WV�^�w�	�|V������u�~���k	�5���
9<t�@@���< u�< t��G�9>�uj �\ j j �߸ ���F��V��Et�}  t�u �q�>> uW�V}[�F��V�^_��  V��3��D��G+G�D�G+G�D^��  V�v�F� �F�  96�u� 3��l�t�Dt�����>� tj j �֋��
 �#�F��V��F�F�t(���6��t&j j �ދѸ	 ����F��V�����
�F����F�  �F��V�^�� V�ȋ��t�d���Lj j �ы޸ ��DuV��j j �޸ ��^�WV�����H��"�^_� WV�����H��"�^_� U��WV���G���G�9Gv��9Gv�N�;Gv�G+����3�^_�� V���L��O�L�O9LsF���O��9Ov6���L��O�L�O9Lv�L���D��G�D�G9Dv�ډG��^�3�^�U��j�^
�F�V�O��t�v�v�FP�i�� U��W�~�t�~��v�v�*  ����W�^�F�V
���F�t�v�v
�v�vP�M_�� U��V�vV�^�F
�V������t�v
�v�FPV�Z^��
  �  V�v�^
�ƍV�������tV�^*��6��F� P�:�^��  �  V�v�^�ƍV������tV�^*��6�� P�=�^�� �  �^�F�V����F�tP�v�F��� �  �^�F�V��r��F�tP�v蝁�� U��j�^�F�V���t	�v�v�'�� U��WV�v����P�>z[���u�>> t��w��S�3��	�vV����^_��  U��V�vV�M����StV��y[^��  U��WV�v�~�Dt���R�d�� V�? j j �ދ׸ ��VW� ^_�� U��WV�v�~�t�V� VW���t�u�^_�� U��j j �^� ����  �  WV�v�~�v�u�@P�������P�E+HHP����Ht!�v�EHP�@P�������P�E+HHP����UB���,�vV�5�^�����P�^��^��vV�EHP�^����P�J�F�EH;�w̋vV�u�5�^�����P�^��'�V�u�EHP�^����P��V�EHP�5�^����P� �V�EHP�EHP�^����P���^_�� U�젶��% ;�u3��6�Fk�
���I�F
���I�F���I�F�V���I���I����% ��� ��
  U��V��9�u3��K�^k�
���I�k6�
���I�Gk6�
���I�Gk6�
���I���I�G�W�~ t����% ��� ^��  U���t� tSPR�v�v�W����3��� U��V�vVjj�	 �t�^�� �
  V�vVj �T��tCV�v�I��D- tHt)HtHt#Ht��D�(�D��P�D�T��P��P� �`�(  ��>F tCjj 褃�u8jj 虃�F� �F�  �F�  +��F��F��^��' �uj ��jj �j����,�~ t�O�3�^�� �  WV���F�  �F����F�  �= t��F�� ���u����>� t����>� t1�6�����V���Vr!��GDu��
�E�U���uNN�ދ�F��}t�}u@�~� t:�^��G�u��;�t�M��v��
���>� t���uj j �
 �V��R��~� t,�}u�^��Gu�E �u�u�E�U�^��&��F��V��F��V�^_���  V�v� �\��9F
u\�|uV�� s
���t�� �v�< u�| t8�L�ɋF��Ѓ���t9t���׋^�w�w�T�^
�( ��� �3�^��  �
  �F�Pj j ����t�~�u�F9F�u�F�Pjj ��� �3���  U��j �~�@�FP蔁�t�F  ��  ��������*� �  V�v�DF�ЋDF�F��V�RP�޸ ����v��v��޸ ����^��  �W��t��t��t��t��t��t3�ø �V���+�;r9Dv9Lw
9Lv� ^�3�^� V�>�0t�t�6�����V��� ^�3�^� V�>� t�6�����V���Vr9tNN����7 ^� WV���t(�����ۉ��V���} t�u�t
������t��^_� �G��G�؃? u����U���� �F����  �  �F
�tHt�� �@  +��@�@� �>( u� �@ ��&�l &�n �F��V��>@ u�@�@�@ �@�@9V�rw9F�r�F��V�+@@��F��V��F��V��>@u� �� 3�9V�r=w9F�r6�@ �F��V��@�@�Ӆj �6(�6�P�6�P�6�P��轅��@  � ��
 �  WV�F
H= w+��.��u���Š۠��!���E�d�|��������v�Du�� �t��m[@P�r[���u� �� �D����D�|�� �v�Du� �t�mr[� �~t� �v�Dt� �ލF���V�F�Pj �DP�J��~�v�DuuV�{ �o�^+ҋG�i�v�F�D�DuVj j �޸ ��E�Vj�g��A�~Ru:�Fu4�><��أ<P�v�"�v�< tj j ��ָ� ���
� �� �3�3�^_��
 �  WV�v�Du�� �D*�����AP�'v�|+|
�|u�t�t
�>�$\�PW��u��6��D
P�D9Du� �3�P����| to�\�? tg��rbS�jl[�F� ;�s��+F���D
�F���D
 �F��E��F��D*�����AP�u�t�F�HPj �F�@@P�Lu�t�v��t�v��u�DtP�D@�F��D�F��D@�F��F�@@�F��6��F�Pj����D�F��D
@�F��F�@�F��D�F��6��F�Pj���^_�� WV�� �Ӌ�����<&u��+�����B�F�< u�ڋ�� ^_� U��F
- r- v�v�v
�v�v�v�H��3����
  �r  WV�~�F�F��F�P�'�u!�u�o'j ����F�V�E�U�= u�"����F��@�F��E#�@�F�P�MQ���}�u�E�	�u�d�E�F�j�5�F�P�u�E
P�v��u�E�Pj W�C���tAV�a�v��F�P����^�����t�>� u�\
�F�V�����t�^����}% t��v��x�F�P�'�~� t�v���F��@�v��	��E�U^_��  U��WV�N
�^��"���?=� u�� v�(��t(,t8��tQ,t0,mtY,Pu� ,s�,w� �� �vW�v�v�v�-��� �>� t�� �vW�v�v�v�� �� ku'�]�p�o�� �vk�]�?uWV�� 9u-u
�6@�6�� 9u)t9u+t� j j 9u)u�� ��� �U�^���tk�E% �d3�3��p��� u3��� ��E�U� ��^�G �E'�})�t6�^�u�E)9G t%j j k��]�~ �j j ku)�]�} �X3����v�v
�v�v�v���^_��
  �  WV�v��-	 tF- u� - u� -� t1-, u� - u� - u� HHu� - u� �v
V��� �~
�}w� �U'��~	u�D9Ew3��F��u�uNk�]�_�G�F�� t�F��t9u'u�k��u�p����qj j �^
�W)�^�x �=��\�v
�|+�tSj j �T+��v
�|-�tAj j �T-�ыv
�V�|' t,Vj���Ku� ��v
�V�DH;D'vVj��Mt�3�P�^_��
  �  WV�~�^��"�?�E%  �E)���E+���E-���u�~
� �F�P�LQ��|�u�D�	�t��|D�F��4�t�F�P�v�DP�v��t�DP�t�t���D�u� �؃uI�Gt��+E� ����E)�\�O��\�G t��+E� ����E+�\�G@t��+E� ����E-��+E� ����\�G kEE;�v�<��v��^
�w�w�^�� ������t&�6B�^
�v��;�s�u�����v���B��~
�E�E'3�^_��
  �
  WV�v�F�  ��� vV�L����t�D���ƉF��^kGG�F��w��9V�vi�ڋw�~� uS�|�tS�\*�\���������t�E�;F�t���t�]���ߊ��*�+F�= �u�DuO�D@t�F� ��D@t��뒋�^kGG;�t'�t�h�\�GHHt
- r- wSj j ��� �3�^_��  �  WV�^kvw�v��9ws���|�E t�v�kww���v��v��~�9v�tj j �\�� ��W�\�G@u	;�v����^_��  U��^�F�G�F�Gj j � � ����  U��WV�v*�D����� t.�Du(�D�΋����@P���DnVj ��~W�\��� P�	�^_��  U��F�� �  WV�~�u'k�E�؉F���F�=
 tv� ,s� ,v
,r,v�w�~u�EH�3��F�9v�tavk��^G���؋F�9u�~ t�]�G�^��_9Gt�~ uǋ]�G�^��_9Gu��Eu��u��~�u
�uj j ���^_�� U��RPV��"�7�D% �F��V��D�T^�� U��SWV�؋v�k��|"�=�}�q�t�| tVR�v�v�v�T^_��  V����k�����"�4�Ë\���@^� U��WV�~�^��"�7VW���j j k��t�X�� � �o�^_��  �  WV�^��"�?kvukFE;�r$j j �\� ��:��u���ދ�+E� �������^_��  U��WV�vj�vV�e���<�u �t�ex��*���E�D�E�D�E�D�|� u��*�+D@��D��*�+D���D�DD^_��  �  V�V�V�F-Ht- t�Y�ڀ?�tR���ڀ�tF�G*�F�^
�����Dt�v
�v�v�v���!�F��؃u	�v
�v���v���� �3�^�� �  WV�~��"�F
=n u�<v�T��t2��ti��u� ��tg,tm,u� ��u� ��u� ,u� ��v�u�� V�f[��u� 3���u�E
  �^�G�����^��G�� �5�bf[�� �^�3��ʋv�F�����Du�96�uVj j ����� �vW�v�v�v�� �E
 �vW��j�j� �ߋF��j ���F	�us�^�N+O
t�G% = �@+ȋE+E;�s�M+MSj �E�~�9Eu� �3�+����؉GP�\�^��F�k��F9Ft� �3��߉G
�F� �,��v�v
�v�v�v��^_��
 �  PSWV���Gt� �Gt� ��^��
 t��9F�u� �3��^��_*��� P�i�^��G+G���v�j j �OQP���u3���މ^��^��_*�^���P�{i�^��G+G�F�;�vSj W��P+~���W��^_�� WV���Du8�D�L�����ۃ�*�؋>��P�+i�t�t
j[�h�t�DHPj]�wh^_� WV���u�D� ��P�_[�D9Dw�DH�DPW�4�_���\�<3���D�D^_� �
 t�G
  ��� WV��3������ǋ����^_� U��WV�~��- t`Hu� - t
- t-� u� -8 tRHu� - tkHHt$HHtnHt- u� �� sq�׋^
�F��t�^
�F��z�jk�u�^
�F�� �th�]�F�^
�����O�3��E�EVPP�)�Ƌ����B�^
�F� �7�^
�F����� �VW�+ �#�^�? t�w �v��׸ �w��	�^
�F�� ^_��
 �  WV�v�~�D�F��M+M;�w+�@�3��DWj �F��~�9Du� �3�+F���+D�DP��ދF��j�^_�� WV�������| u�| u3�^_��L�ǋ��@��Wj �L�t�N� ^_�WV�����W��DD;Ds%�E+EH;DvWj �D�t��^_��D�ǋ����^_�U��PSV���^��GG��;Gs(+w��V��@PQ��_���^�� t�O�^��F���^���  RPSV�
 t����^��GH;Gv[�GG�F��>< u9Gu�G�7�_�  �>< t�^��G+F�P�F�P@P�i_���^��F���v�� �^��F��:�� ^��3�^�� U��V�N
��- t- tfHHtp� �vQ�v�v�v��^� tA�Gu;*�G�O�����ۃ�؋6�� P��e�vj j �^�wj�����vj �J�3���9�v�v�v����^�? t�w �v�� �V�8��v�v
�v�v�v��^��
  �  WV�v�|"�~��F
=~ u� v���t/,t2,t@,tH��u�� ��tz,u� ��u� ,nu�� �� �  �� �DuV�5�� 3���� V�v�v�m���< t�t� �~��- t- t�t �v�� ���}�� j j ��T �x ��j ��d�v�dV�5�s�uq����V���^��t03����V�^��'��7�f �\
�F�V�X��tj j ��T �x ���vj hV�^�w��\��@P�l�j�[d�^�O�S�^��7� �v�v
�v�v�v��^_��
  �  WV�v�< u�\��*��>���%��_*��>����_*��	�\��*�2	��2��F��| u3���t�hZ[�F��D+D��- ;F�s�E��F��FtY�> uR�\*���GP�cVj jj �E�P���| tVj j�t�v��t�F�P�ncVj j j �=�Vjj j W��� �\*���P�GcVj j j �E�P���D�tVj j j��Vj �E�Pj���| tVj j�t�v���F�P�c�> u)Vjj j ���Vj �E�Pj܋���Vjjj�W��Vj�^�^_�� �  WV�v�|"�F
=� u�Xv���t2,tM,te,tm��u� ��u� ,u� ��u� ,pu��W�|u3��� ��D�t7�L ��8V�v
�v�v�v���V�5�;3���.V�v�v�����t��~��-  t�< tO�t �v�� ������ Vj j �u��� Vj j��j��a�� j ���u���D�V��5� �~����u� 3��)�^��'��\
�F�V���tA�|u�^��u3j j �^��% = ��ډV��޸� �)�< tj �v���T �x ��V�@�% = �@���߉~��% = �҃� �~ t��^	W��'��^��!W�v�^��7� �v�v
�v�v�v��^_��
  U��WV�v�Due�~��% = �ۃ��D*�؋ǋ>��	Q����`Vj j �߃�����j���\*��>��P�`�| tVj j�tj���Vj�#�^_��  �  WV�~
�v��"��=� u�+v�h��t,tL,tQ��t^,tI,�u� �J�^�G+GHH�D�L
�D��D�D�D  �D �d
��O�3�3��&�vV�%���vW�v�vV�m�� �D
u�� V�t�*��9Ds�|�D
$<u�^�? tj W�W ��� �q�d
�3��&�� �~�F��u� ;�w���V�E�P�@�D9Ds�D�D+<�߉|�D9Dv�v�V�D+DP�;Ds
Vj����vh� �vj j ����vV�\ �B�v��~VW�C�^����G�;Gw�v�9w	�G+G�F��F��w�G�vSV� � ����v�v
�v�v�v�z�^_��
 �
  WV�v�Duq�~�\*��D�΋6��R���N���^�^��F�����v��F�Pj��Q�#��v�j j j�{��v��F�HP�F�HPj�iދE@�F��EF��F��v��F�PjۊP���^_�� �  WV�^�~�w�Eu9vu� s� �3��F��]*���Q�3^�F�  �F� �~� t�F��ƉF�@�F�~� t����F�F�@�F�+F�F��^;Gv	�GF�F�W�F�P�~��$+�P�EP�HދF��^9GsF��	�GF�GF�W�F�P�~��$��P�EP��^_��  �  WV�~3��F��F��E
% �F��^�F+ҋ�+w�F+G�F��~
t� �~�uM�E@;�tB�t>�E@;�v6�~��~0�~�}*�E�F�@;�s"+6@�u��E;Er)�E+E�E��V��� +u��6@;us)u��E  W�u���9Es�u�vW�v��i��F�� �V��v�� ���u�u9N�t�~�u�� �F�� �o�V��E+�=��u�u�t��uU� �F�� �K�EE;�s�u�t��u4� �F�� �*9ur�u�t��u� �F�� ��u
� +u�6@�E
��2�% 1E
�t�^��~� t�^�? tj �v��W ��F���^_��
 U��WV�~�v�= u3��
�U�����g���EH;�s�uN��^_�� U��WV�~�v�= u3��
��]���g���H;�s�5N��^_�� �  WV�v
�~��"��Hu� Hu�� Hu� - u�Hu�&Hu�:- u�:Hu�- u�Hu��-y u��Hu�Hu�(Hu�'Hu�Hu�Hu�Hu�Hu�Hu��- u��Hu�Hu�Hu�$- s�3- w��(�  �^�G�u)�~ u� ��v���tV�?V[��u� 3���u3��E
�E�E�E�E�^�G+G�E3��׃= te�5��U[���vV�v�v�v����vj ���ԃ>� u;�vW�v�v�v���vV�u
j�M�j�<Z�} t�j �.Z�m�} u�d�v�D9FsVWhHj j �e���@�D9FrVWhP��\�F�V���t��D@u׃>� uЋ��.��5��9Ft�3�����v96�u�\�F�V�x��t�D@t���F+D�E
9Ew�EH�E
V���v�EE
j P��T �� �	���v��vjj j j ���vjj j �v�����u�vjjj j ����+���F�E�v9EsVW�Vj �T�v�U�E �v���u@�]]�F9Ew	;�s�u�);�u�uF�9Ev3���EF;Ew�v��u+u�F+ƉE
�u�vj�0�v�u��v�� �E�h��EE
�_��ߋF�Z�T��^�GtW�v�)����u�~�����~��F���.�^���+?�v�W�v�v�z���^�3��G
�G�v�w��^��G9Gw����vS�����v3��EP�P�v�} t�M��EE;Es�E�vVj�lV�u�C�%�vWhIj j ���vWhQ���F�E�vj�>�v�v
�v�v�v�"�^_��
 �  V�F-	 t- t
- t-� u�-8 tlHttHu� HHtHHu�HHu� Hu�� Hu� �~ r�b�^
�GG
�F�� u�N��vS�v�v��c=��u�Q�vh� j�j P�u��@�v
3��D
��v
�DD
u�� �| u�^�G@u�� �|
 u�L�� �L
�� �v
�| u�D
  �� �D9Dw�D  � )D� �^�G@t�v
� �v
�D9Dv�D+D�D�DH�D
� �D��v
�DD
@;Dso�| u	�^�G@t`�^�G@t�DD;DsL�D�G�D
@;Ds��D
�9�v
�DD;Dr�^�G@u�D+D됋DD�DD;Dr	�D+D�D�vj�z�v�t�O��^�? t�v�v� ��V�p�^��
  �  WV�v
�< u� � �D+D�F;Fs�D��P�4��c���t؋^
��G�F�^
9Gv�G+FP���FPNNQ�sN���^
�FG�G�N����,��*��y�*�P�v�EP�AN��3�^_�� V9Gv�? t�7���	�*�@@�J�u��^�3�^�U��WV�v�D�t�4h� �t j �v��W��v�~�D�E
�]�*�E^_�� �  WV�v�F
�F��D�F�~�F�9Ew�F�  �v
�ߋF��l�P�F�P���~� t�^�*�&�P��K[�N*�Q�F���K[9F�t�F��F�;�t���u�3�먋F�����^_�� U��WV�^�? u3��/3��7��v�DP��a���G�*�@@��^9wދ^��+^_�� U��WV�v�| u�LV����Du�tj �lՃ| t�~�u�u�\�U�� �c�^_��  U��V�v�d��| t
�t�1�V��^�� U��W�~�} tj j �]�� �V��_�� �  WV�v�|"�= u	�D�u�6�} u��D+DH�F��E�����F��E;Ev�E�F��E�F�v�~ t�D@u�E �EE
j P�T ��� �։~��Dt�� 3҉V���9~�v�~�F��F�^�9
u� t�F� ��~�� �F�  �D t�4h� �t �F�j P��W�XVP�F�P���D*�~��ۃ����P�RVWj j �O�VWj�v��v��v��eҋF�9F�sVW�F�@Pj �F�+F�P���D�u�^�*�@@F�G�F��F�96�u	V�u
j�<�^_�� �  WV�v��r	�~�u����u�>> t����C�> �>@�F�@�v�v�v
�vk���@��@�wh4�w���p� �>  �>@^_��  �F  WV�~ u�v�]��F�F�j/h��F�P��J��kFP�M[���u�>> u�H��I�~�3��~��jh�k��P�J��F9vw�j �v��F�P�N�Q��F��F��~�s�F� �F�V�F͉VϋF�F��F�  �F�F��F�  �@�F�3��v��~�� ��ދ�^
���k�߉O�G  �ˋڋ�^��ىW�G  �^؋�� P�^�X�ىW�w�F��^��\�F�j&P�}H��= �% @@�v��F��G[F��^��N�ىF��^��G�F�- �G�^��Gt�v�F9vv�Z��~��v�T��;V�v�Vȃ>> t�F�P�nQ=v����o��HtHt#Ht�D�F�+F�^���G�4�F�+F�^���G�F�+ǍL+���^�H�G�Fȋ��+B�+Gk��@�F�Pj �v��ۋ��~��It�v��K[��^_�� �  WV�v
�t�\*��>��P�O3��F��F��v�=hDV�G�����F��~
 t�v
�v��^�+���PVW�R��9F�s�F���<
uF�< u��~
 u�^�F���^�F��^_��  �  WV�~�]"�F
�7- t-u t-�KW�v
�v�v�v�9ۋE+E�F�W�tj �F�P�5�3���0�F9D-tk��|�A�D�D  �D% ��W�v
�v�v�v���^_��
 �>@ tj jj j h@�@� U��F�@�N�V�@�@j j j j h@��3��� �  ��*�F����F�@�F�3��F�Ph�ɍN�QPjPPh� P�v�Dɣ�= �% ��  U��WV�F
Ht0HHu� -�tDHtJHt\HHt�v�v
�v�v�v�m�� �v�]�F�r@jPj h@�YG���n@ �@  �ƋF�r@� �v�D����p@�D����v���D�p@�jQh@�DP��F���OV�D[����Pr�P �6@j h@��F��WVh@�F���>@�^�_*��6�� P�FM�vj j h@jP�5�3��^_��
 U��V�~ u
�v�.Y����v�>� t�u�hj j �֋�����^�� U��>� tj j �����V����  U��>� tj j �����V�_���  U��>� tj j �����V�?���  �  V�v3��D���F��F��F� ��*�N�V� jh~͍F�Pj jj j jj V�j�^��  U��WV�~�u�$�u�t�FX�D���׉D�t�t�����kEE;�w�^_�� U��V�v�u	��3������F�t@�޸ ��Vj�x͉6�^��  U��F�t@��  �  WV�V����"�?�ڋG= u� v� ,t,tb� ���tHtHt	� �� 3ۃ�+r� ����*�+D= �tC��W���w�Y�E=��tfW�6��g �6�Wjj j �)� �M�>�u� ��>� t�W�6��9 �}�u�E  �6�W�"���E�t���>� u�� �M@��3�^_��  U��>�s)�� �^�O@�F��hv@�����9�t�6������  V����"�7�>� tA�d�D���6�V��>�r#��  ��� t�w���6���hv@����  ^��  WV�^��"�F
�7=e u�v���tQ��t[��tr,u� ��u� ��u� ,u�� ��u�� ��u�N,u�,u���u�,Eu���F�^��"���t�j j �֋t@�g �k���v�v
�v�v�v�2��vV�3����d��>� u��vV�v�v�v�n�݉v�V�v���G�>�t�=�t�F�^9Gu�*���$�^9�t&�����j j ��� ������~W�k��D t���L �t�d����v�WV�v�v��F�9Du"�} u
�L�v��� j j �]�d �������v��t�L�v��} u� �u�Q�� �D u��d�3��σ|�u�����t�Dt�~WVjj j �l�d��M�ىv����G u�=�~�]
�F�V�8��tiW�v��v�v���F��^�9Gu��t�} t�u��ŋ^��O�^��F��G�Gt�~��tW�v���W�v���~
et�� �^��O�� �} t,�]��
�F�V���t�^��g��v�v�]� �V����^��u0���
�F�V���t�^��g��G��WS��v�v��e �^���tN�G��WS�B�Dt?�6����v��ċ���"�7��O@�do�6����u�L��F�D�vV�D�v�v
�v�v�v��^_��
 �  WV�v
�u� �V��- tQ- u�� - u�"- t<- u�MHHu�g- t(�v
R���F�=��u��^
�G�vSjj j ����~�D�F��d�WV��} uWV�s�u�e�} u���j j �tk^��P�t@�( ���A�vj j �\�d �����t�'�V��- t&- t'- tn- u� - tIHHtE- u� �I��|�u�d��� �ދG�F��wk��8� t�� �F��Ǩu8j j �^
�w�k��~�5W�n�j j �޸ �V�a��|�tk|�\�y
�u� �� k|�\�q
��`�� �vV��p�D�L�u�DH�Dk\\�?�u���D�D9Du�D  k\\�?�u��vV�a�D�t�Ǩtj j �^� � �����9Ft�v�c�^_��
  �  WV�~�M�kuu��t3��� ��u� �� �F� �u��t�{;[@@F���kEE;�w�ku�]�x�eǋ��@��E��j j �׋t@�f �K��F�  �u�~��u�t�%;[��;~�v�F����^kGG;�wكF��F�F�@@��*�;�v��*�+F�HH�F��F��F�F��F��^�G�F��v�DF�@@�F�jh~͍F�PSjj j jj V�*�= �@^_�� U��WV�~��� w
���t�� �^�w�~�^kGG;�vZ�|� t>�\\�������t�ȃ� ���;�t$���t�ȃ� ��ȋ�*䊇�+�= �t��먋^��+G� �������^_�� �  WV�^�t�F� �^
�F+G��F�  �^
�F+G�F��^�w�^kGG;�v<�t�t��9[��GG�� �F��9F�r9~�r�~����Ƌ^��+G� �������^_�� �  WV�v�>�u�|�u;hv@����% = �@�F��F�  = ��% �F��^�G+G�F��|�u+3��.kDD�؋��u�� t�k|�\j �q�J��kDD�F�D�����J�tG�]*���P�MB�EF��F�P�E
@PjċE+E
HHP��A�v��u
j��A�v��EHPj��|A�� 9v�u�E�F�j �BW�v��F�@P����% = ��$E�F��^�*���P��AW�v��v��% = �$P���t�M8[�F�W�v��F�@P�t�v���W�v��F�F�@Pj �~� t� ��F�+F�HP����uG�^�G@t>�F�9Ds69v�u� �� �E*����P�EAW�v��DF�@P�\\�P���~� t
�F�@@F���F����^kGG;�v��^_��  �  WV�V��- r- v�@ ��  �V��v��4�~u�� u�@ �$�F  ��~u�� t�W�= u4�F��F�v��v
�F�P�v�DIP�v
�}���u��F�^% ����� ^_��  �  WV�v�~VW�@IPV�H�tP�= t� ^_�� �  WVh��;[���u� �@�~WV�6��V�v�-IPV��F��tP�p= t��VW�f6���~��� V�Y;[��^_�� U���v�
IP�v���� �  WV�v�~�v�v
�vV�F�P�<I�F��t�F���
9v�t�F� �v��v��F��tP��= t�� ^_��  �  WV�v
�~V�v�vW�F�P��H�F��u 9~�tj�F�+������RPV�L���F� �v��v��F��tP�= t�� ^_��
 �  WV�v�~VW�v��HPV�� �t= t= tP�Q= tܸ ^_��  �  WV�v�~V��HPW� �t= tP� = t� ^_�� U��V�vV��GPV� ^��  �  WV�v�~WV��GPV�n �tP�� = t� ^_�� U��WV3��~��DP��EHHt	��������� F��r���E�tHt�2��E����E= ���� 3�^_��  U��WV�~�>��t�>���� �����u3��M�V�t
Rh�A�G4����� w#3ۉ~��s�ǋ��8��tC���*䊇��Wh�hjh�B�:��� ^_�� �  WV�v3��th����ta9>�t	V���tTh�Bh�A�ƙRV�� �P�� ��
9>tWjP�� �h�P���*�P�����"���jQ�GIP�3H�� �P�+Hhn�%H��^_��  �  WV�vV�3[��;~sV�v� �|:u��Ph�hr�v�| ��FF�hz�v�@3�����9~w�v�h��DP��4��@�+��< u�< t
�~VW��2�,�~W�53[��+v�ލL�Q�v��P��5��h�~��W��2��^_��  �  WV�v�~�u�F�	�v�cHF�F��F
�F�� �?%t�F���F� �F��^��?.u!�F��F�P�53[��h��v��4��F��F���B �^��F���=u tLwW,%t,+t,t,t(�E�%F� �<V�^��F��7W���,�^��F����݋^��F��7V�2���V�^��F��7��FV�22[��^��? t�H�� ��+F^_��    �                      MS Run-Time Library - Copyright (c) 1992, Microsoft Corp     x ������������������������������������
���
�
����������������������    ��      F   �2 �S &O �N �S ^S 6Z d[ �V .X fT �T fV �V \O �O (P �P �P Q �] V\  �\ �y  z �}	 N pN �N 6Q �=  �A  �= *@ �@ ��  �M �8 �8 P9 n9 � ڄ �2 �2 Y 0Y LY �Y   ����             �       �  �     �   ��� � � ����� ����� � � ��� � � � ������������������������������������������������ 	
     % '  '   ! " '   '  ' ' '  
  '  	 '   '  ' ".<@HN\bj��   H P K M S  	  
 	   G O �   �   Q I v � t s u w ;, = @' B c% a& e(  0      	           � x1 y2 z3 {4 |5 }6 ~7 8 �9     -  $             .  . F    A    Y /  / S    D            �  � e     �  � f     � ! � h     � " � i     �   � g          ��    � # � j          ��    �   � k   	 �      �  � p     �  � q     �  � r     �  � s          �  � y     �  � z     �  � {    N      � % � �     � ( � �     � & � �          ��    � 1 � �     � 2 � �     � 3 � �     � 4 � �     � 5 � �     � 6 � �     � 7 � �     � 8 � �     � 9 � �    z      ) � �     * � �          , � �     + � �    >     � � ��   � F� ��   � r� ��   � � ��   � 6� ��   � V� ��  ^   �����    
�   @       P����    
      !        ����    
�           ����    
�           b����    Z             b����    ^      $       b����    _      D       ����    �       �     {                �����    
�   @       P����    
      !        �����    
�   @       P����    
      !        ����    
�           ����    
�           b����    �           b����    �           b����    ^      $       b����    _      D      ����    �      
 �     {                �����    
�   @       b����    �           b����    �           b����    ^      $      �����    �       �     {   ��            ����'    
'   @       P���(    
      !      ����)    
      @        ����*    
*   @      
 D���+    
      !���     ����,    
,   @      
 D���-    
      !��     ���.    
.           ���/    
/           ����0    
0   @       P���1    
      !       b���2    Z             b���3    ^      $       b���4    _      D      �B��&    &      v     {                ����Y    
Y   @       P���Z    
      !      ����[    
      @        ����\    
\   @      
 D���]    
      !���     ����^    
^   @      
 D���_    
      !��     b���`    Z             b���a    ^      $       b���b    _      D      �B��X    X     
  
     {                �����    
�   @       ����    
�    $       ����    
�    D       b����    Z             b����    ^      $       b����    _      D      x����    �       ^     {                �����    
�   @      
 D����    
      !���     �����    
�   @      
 D����    
      !���     �����    
�   @      
 D����    
      !���     �����    &�   @       b����    �           b����    Z             b����    ^      $       b����    _      D       4����    �       0     {   	             ����!    
!   @       P���"    
      !       ����#    
#   @       ���$    
$    $       ���%    
%           ���&    
&           ���'    
'           ���(    
(    D       b���)    Z             b���*    ^      $       b���+    _      D       N���             �     {   
            
 D����    
      ��       b����    Z      4      �3���              �     �   ��           � &                         #  #  #  ����EDIT.INI  EDIT.HLP  TEMP  TMP  	   	,.;:(){}<>[]"'\/~!@$%^&*-=+?| LPT1  LPT2  LPT3  COM1  COM2         �����߳�������ߋ�߲�������                                               d     �                           _C_FILE_INFO=                                ���                     ��            ��PX   	��            (((((                  H����������������������  � � � 	 �� @    GHIKMOPQRS  @ l @      �  � �  �����������������߼߷������ � * ����� �  ����� �  ����� �  �� �       
      
   , . - :  �$A �    ENU �  ��xyz{|}~�       0. !"#$%&21/-,    ��2 �  �            ^�P�b�L���    ��& �  ���    P      P   �  @   t  �ĳ�ڿ��� ��ڿ��. �  �� X\`d � 	 �        
 �  ���  �      �  � �  �0 @    @                  Z ^ [ \ ] _   " . (   " .d f h j d e g i pqpp��ppx��� ��ppxp    ppppppppxppxp    �� �  ���'$���	�
��������    ERROR 255: Unable to load string resources!
  *.* 
 % %c: %s\ , *?    [ ] [X] ( ) ()   %u  

  %c:\... \...  \ ... 0123456789      ���� �  �<<NMSG>>  R6000
- stack overflow
  R6003
- integer divide by 0
 	 R6009
- not enough space for environment
 � 
 � run-time error   R6002
- floating-point support not loaded
  R6001
- null pointer assignment
 � �� ���    n <0RB��� �  ��� ��O����P�4 PˌÌ�H�؎�� � ���G����H��� ��������+�s��+�����ڋ������+�s��+�����¬��N���F��$�<�u���<�um�¨t��2� �3ҭ�����Î�������t&��� �t�� �܌�@����&H����Ë> �6
 � - �؎��  ��֋����.�/�@� � �ʎں�!��L�!Packed file is corrupt �DSC$�`��0|�4E�                              rt
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              A<�R                                                                ' ppppppppxppxp                        Aqpp��ppx��� ��ppxp                        |�D�D X� �tA� W &��&+�&
�- �.�ﱸJ3��/.9�w�� �w.�ﱸJ�/���t� ]^_ZY[X�  W� �.�ﱎp�_� �+����������+��/ �p��&��� �> ���6 �|�D���I u��&�^�&�s�@&�Z�H� ��&�t�&�v�Ì�&�֧� ��&��&��ۥ�� &���&������˜X �P��X� ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �X                                                                                                                                                                                                                                                                                                                                
-- More -- Line number:                   u    A          =t=Kt
��Ht.�._�.�_.�e.�g�c�<u�ڀ?���u��� 3��
�u����PSQRVWU�.�.��,u_�b�'�(�t���6(Ƅ'�'�r(�>�(���t�>�'�(G&�G���O�,�>&�E �=�>GG�� I�,u�� �6�
�t3<t(<$u�
�t&<t<*tM<1r<9vu���ج
�t<u��6�� �&,�6�(��<��u�,�6�(W�� _� V�6�(�tK�< t�<	t�NC�tK�<t	��2��^�^�i�V�6�(,0���t�K�<t�< t�<	t���t�t�K�< t�<	t�<t���CN�t�K�< t�<	t�<t������릋6�(�tK�<t������6�(�u�&,����ϋ>+σ�&�M]_^ZY[XË6�0 �!�6Q�B Yr�G)(�>�,����<ar<zw$_�3ɬ<t< t<	t<=t<tA��Nì�����I&�>&;>	s-W�u�VQ������Y^u&�= _tQ&�	+�2���Y�������Ë6�t.;6t$�&���2���t;6t�6��;6t��6���6�t� r� r
�
�u�F�� �6��;6�t;6u�6N��V3ɋ6�t";6tWS3�� �	�
�t
�C���6���[_^�WVQA�>;>ۡ+�;�����t�+��>���;>��Ӏ�t���r#W2��+��t�>�+����Q �6_�E� �>�>Y^_Ë6�& �t��KI�t�$_<Ar<Zw2E�$_t�Ë6�׋+�s�+��;6u�6ô���2��>���#�ô�>���6 �!�" À>" t��>�*6"�6 ��>�6 �!��ô��<	t� < s
<t<t��ù".*�2��Q��Y�!2�+�s
� s��!���VQ��Q<	t&< s<t<
t<t<t�Ȱ^�� ��@� XY^ð � �����û ��6;6v�+��
 �6�+��_P�ǀtI��
�t:�t��3��6B�uQV�D�_ ^�;YC�2 ���9 �:�g�� ;6u�>�Z���t� C�
�u�π��C�X�ð�:��
�5�
 3�.�6��Rt���X0�����
�u�ô���!2�<t2�&��:&r&SQ��>�Y[��:u���!�
��!2��"�&��1 �(  �*  �&,�3��؀&���> t�8�h� ���6�'F���2��v� &�%��<t���&)%�
�@		
_@	0	qnCBAtswu@?>=<;SROGPHKMIQQ@	A	A	~	c	���	�	��	~	�
�	�
m�
4
*
F
q
?��
X��� ���� u	��� �������'P�t X����#��XÃ> t�P���X<It	������>* t�*�6*���2���Ë6*;6(r
;6%t�(��'������*���u�Ë6*;6(t���������u�ù Q�,��[�>*)(r;>(v�>(�1;6%s��'��'FG��>%Q�����X+������>* t�P��6(N;6*u��6(�������6*�q�Y��t�6*�6%�6(����6*�tJ��'�t�6*�t9N��'�pt/�����6*;6%t ��'�Xt��������t�6*��'�At���I�� t"�6*;6%tF;6%t8�'u�V��^;6*w����� t��6*;6%t�F;6%t�8�'u�+6*������������  øD� ��2�!r�>8t�@ �ؠ� 
�u�2�B�B�(��&�����6V�6;6u�6�6^;6tV� ��'�*���t^;6u��^�6*�� �X�*+��Q���Y��Ã> u-Á�-v5N� �.!Q� �U�� �o�� �J�Y� �.!�� ����Q�7��-����u�<t^<t<t�<0r�<9w��2sވF�'��֋ξ-+�3��5�&��ج,02����ء��˃�vQ���Y�;t����%�2�P�6�k�X*2���X<u*á�	��@�����&,����6%�.����%�&,�ÿ'���(�%�*  Q�)�*�������ۃ>( t���w��̀6,�2,�Q�#t��w2��	�Y3��؀&.�,t��À,�,uj�6*��sj�6*��'���6*���*��F�6*;6(v�(;6%v�%
�t�P�\�X�6*;6(tP��'�����X�����F*�u☋�� �6(��r����6%��tF�6%;6*tN��'��(�'�(������*���� ���  �6*;6(s(���F�����6*;6(s��'�P����F��< t<	��(���/��!
�t��!��
�u��!� �Q��Y�� ~� ������  /REINSTALL /BUFSIZE /HISTORY /H /MACROS /M /? /INSERT /OVERSTRIKE  �0�!=t����� ��B�tt�E�t\�M�t\��}tD�+�utm�4�mte�7�etf�?�]t^�"�Uu_�E<=t�c�:�U�Y.���.���.�� �.��@끻��C
�t
S�д�![�� �(.���_�.���V�.��u� H�/= Ht� V�Y=s������;�v��P�, �I�!���	����[ã�ȣs�w�}��{�+����ˎ�&�� &�� �_�a�.��^� =���u
��t���h.�� t&��.��@t&� �!�������<=u8���� �F �Wr+.��t2��Q����.��t2������ ��������u�L�!��'WS��u�GKu�[_VQWS� [_Y^�=��� &�&+	+�vP� Xr"&VQ����&�>	�2��Y^�2��&�>	��WV���<t@<$u9�<t7<$t<*t<1r<9w&�$G����|<Bt�<<Lt�><Gt�<Tu��Ī뻋�^_+�Ë������rW&�	+�2����_&�&�>	�QVW�>+>+�r|��rv�;sy++�vi�6+�;6v�ϋ�OAP2��XuO�>�6�>��+NO����;u�6�6;u�6�;u3���_^YË6�6�;v��>���6�+���ON��GF��>�6;6v���O�+�2��>끴	�!���	�!�F�<	t�< t�N�V&�= t	���t�^�X�3۬,0<
s�����ۘ���N�2��6;6	t����=���� ;6	t�����
�tشb<|t�g<>t�l<<t�t<t<$u���P�$��X������An incompatible DOSKey is already installed.$Cannot change BUFSIZE.$Invalid macro definition.$Edits command lines, recalls MS-DOS commands, and creates macros.

DOSKEY [/REINSTALL] [/BUFSIZE=size] [/MACROS] [/HISTORY]
  [/INSERT | /OVERSTRIKE] [macroname=[text]]

  /REINSTALL    Installs a new copy of Doskey.
  /BUFSIZE=size Sets size of command history buffer.
  /MACROS       Displays all Doskey macros.
  /HISTORY      Displays all commands stored in memory.
  /INSERT       Specifies that new text you type is inserted in old text.
  /OVERSTRIKE   Specifies that new text overwrites old text.
  macroname     Specifies a name for a macro you create.
  text          Specifies commands you want to record.

UP and DOWN ARROWS recall commands; ESC clears command line; F7 displays
command history; ALT+F7 clears command history; F8 searches command
history; F9 selects a command by number; ALT+F10 clears macro definitions.

The following are some special codes in Doskey macro definitions:
$T     Command separator.  Allows multiple commands in a macro.
$1-$9  Batch parameters.  Equivalent to %1-%9 in batch programs.
$*     Symbol replaced by everything following macro name on command line.
 Insufficent memory to store macro. Use the DOSKEY command with the /BUFSIZE
switch to increase available memory.$ Incorrect DOS version$
$na /P:1e8,12
rem DEVICE=cd1.SYS /D:banana /P:1e8,11
rem DEVICE=cd1.SYS /D:banana /P:168,10
rem DEVICE=cd1.SYS /D:banana /P:168,9

LASTDRIVE=Z
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       ��\� 0;�si��-D�%������ ��~��ر����S3�S�PKLITE Copr. 1992 PKWARE Inc. All Rights ReservedNot enough memory$� 	�a�!� ����OO����������FF� ��� �2�����;����<����A����c����d����e����f���r���Jt�s�3�3���Jt�����Jt��Ӆ�t��Jt��Ӏ�r��Ju�����.����
t:3ۃ�t&��Jt�r��Jt�����Jt�����Jt��Ӏ�s.��,���V��+��^눬Ȁ� <�u��3��Ju����Ӏ�r���Ju����Ӏ�r���Ju����Ӂ�� ���3�� S�؋ȋЋ����� 
      	          	
�  �
Copyright  (C) 1987-90  ( Central Poi	   Software, Inc. �� � ���
?!�CN�Q:8D�cur0rt_.fil�`4� � &�I����  ���,�'������  �3�S��4� \ �>�   �G� �9�ˀ�r	� (?��u�W�3�E P�!��r����0  �ģn= s
�?&�  ��`	3��l��� T�6� � r��V&t0�>(JQ.x.�.2	PR
�+��
(
)��

X

�
	�/� �t>��wu��.�  t	�2��?��ht����ij$u� ( ������� <7��Ȣ@A�J 
�Er���-���P��uhIua� �B����/��_9�P;�<k<<88<t4�u,�O3  Ҹ02�Q�Y��v� � ��ѹ0(	���	��
 C��$���*�!� ي�p���Ʊ��  ����	���6'�Yb�����6�.���u ��s��f'� ���%
u� ��>nr�4� qC�	Der�� �(�u��o2�H<�u��A	AJ�ݍw �A� �.G �,r��G�.

� M�ܰ�B�jI"r)��=v��  �K�f@=��s� ��ӜB]  �uر��3�����。���  �&Cr��6 #�o�b�D� @JI�d2&� ,L�h�<((���_�<
�r(
��[&�(6erun�: �; r�Q �j���<+�3�����3��ӫBKu����?Pi��-� (��o=r	�?=(@�n��Ѡ�R����� kM���~s<uP 
�n�$<?t���
��>?u�o�T �y���S��F�DIF�(nO�J LH
2r��s���  E�6����j�u�3 @ uC���� t�P[Mf�� �W���&3
�h�;uh�;@t�5GGC��߁ �X��3�����b�&͓�ܡ�Q�����s���A�mm�B� m��d�>���~��>���b�I=|rS "�~��'�Đ
@ut�� &�	�����(����  & (�U&�PW�}�$ (�� ��_X�u; (&�]�u$  �M&Mu�u%�� �r;Mw�v0"u+iF�	e%[u �TxK*D�;Ae�6�ׇ_+t��J�VB��6t�� ;���W�����_W�)P�_8�
 � -�t �Pr���r�;U@t�>>��Wz�v`3��I�B�_����uA�t3�/��fI����E‬Et���B���	�� &�-��P� ⵡ0!t&$@���(����
�
��:��>t�!�)�^���^z�p�f��P��s'  +�7�r�t�<Yt<@)Nt<Qu��A 
��� �G�� 0=��t.�����Ha8���>�H�Z�]Ls	*�'�C�*�GX��)���=�H�t����=P �t
=�t=��u
	&;�u���&�}�:(�.�: ���!�>r@�t(�d�Bj����0���Uu�v�c�����(�(�[��'�pӀu_ �*�1�uM
�P
����GJ�c'���c �S0(>󫣂� �L��H�����  2��O�)r ��;r{&��s����u���$&�U�UuJ�bt�	��� _钋� �G 
 @���.B�8ƚ�#�*sE+�x����@9�Ȓ����G� l��� !�J 6�.�|�\�\�(�=�_�P0t	U�v�'P1��%N&�&6�1����r(�e�E�	5�`*��	���i�����8 ��:  ; ��k�P<ds��x������<Ttʞ�{ �@�k��U)��b����a��&� �:�U��������}�-~�/* �:����M'�C�-��;���)�4�b5�3��c�b+\7�7T��W�>j8�M��٠H�HϖN5� ��U r�(H�.<�w�l���A����  ��!�� �R��WSQ�!RVWU��RY���ł ��6������᠔nt����K�^@0Wu	�6�'V�&� X6�	%Y^��s�F�@�t:�ȣ> �68 ����:@< .�3ۊ$�<�T\:�t�@ u��@М' @�,���]_^ZY[�PR"wM;�r- ��K$�� ۉWZX� �S;�tP��8FTD�U����x�����Av �r
U
0%��EA��!��rU-�}w�S P���r
��X�� �À���N������� ��r��&��P�QVW�.�&a)�ܐ�p��6' $��.rv��@ ��_^Y�PW
 o��;�r�>@�>��V%�� _�U����?3�p�u �� ��
 J��tz� �
%�u�@b�� �GD��?.t*� �-�< rG�w@d ��t@��	(>6<�t;�b -���45u"�G
 3�t� <.u;٪�u�� �		
s���(�e��t�8� �t
�O�.;f��[�Q<~w  <ar<zr�;���  2��Y�:���."/\[ A]:|<>+=;,��
���3ҋ��������0\�uAe=��	�v3
�� ��
&����!A��t&6�
��*ĸ�H�@��d ��������
@�p����t �N��hr���&�OON%�:\=� ;�u�XB�p��ZCG�Iem�K5R
3FF��P
�7GG&�5G�`�w�O �����ȋ�@��+�v��QB'R�ߋ  J+�rA��KC�y}�;������BJσ�C:��_3ҋ��)�0<�`A����t% T=��u��
t�/�����@�@��؋�4Ċ���u�
I�PBDB��(=����9��OPV�|H �2x�tG�)JB����?	���pŘ���뺺�IqMT�P���v���Q ��\(�ú�����{��u��,JD,�@�@1��u� @V�6�����XYu����u%�� R;�s�) #&�nt�?�2��}`%	 h%r�����"T�sۉ�Ĭ�7R���k�s�"��DG�1B�Z��IQ2"��";A��u���$}.tD!��r�ރ�e;�$��C��WU���=u7�΃��	�� s*��UE�B3Ǉ �;��v���\�t��hb��`�>L�Pe*�B �P�Ӎ  �G�\�~�^��>�H��t �3������%HB�  �b��r�q�`�9������W�EϪ�wq�s3�� ���!��* � ��	+Ȱ\�}�:��E%���_�WdW ��e��U P����l ���(� ;@"�tC�d��uBA�����`b�����_��4PX>Eu���Q�jIF���-S�&�2�
5��,����Ж�����Q3�;�ZYã�  �Yc+�@
���r(��A�ø#�@�z���$�Q� "z�G(nu����5�0��*
�t(^�~ؠ~uCB�y�6�"�C*�0BJ��%UL!������NF\H&� ӗ]�`��x:\ �J�/TEST  �/PARTN��)/J �YU��59P��Lt&#�  '�'�'�'	((  ,(6(E(	W(
n(3a(z(�� lzSav SUBDIR;mVE�MPXRO[6.M s ked partions='D�A :\&SAV.FI��L��0Eq��L��.�8��  �L/�,�r/tJ <Ar�<Zw�,A� ش�!���ӴP��X:�
�u������Yn[��H��a�,dC� =-�  6r���23ҹ 
��?�r�;�uǎ��3��h�T�r�?�R��u�u0��&�G	< 15|�&�v+�9umw딍>�!33�"R��,�@��G"��3	�< u�&��G2(4�؈G
� ��RT��	.-����5�-� R��
W,��E+:�*E��� �0�(	�$��
� ��g��l��Pe7��l���@�z���E��;����Ơ����� (�����2$������Pt����:��4 r��<�j\Q�\�/�(��/�3Dy1�\#S�G16��,� 2�A��r 9t-<Qt)�>#=l�<Au���$,0v�:w�H����"�5���( v���r�u쐴
��!$��8 ʋ>���$��t%� @=70���5
P����㋿b��`���A��#���Ba� ���@ �!$/�����雷�R�ѥJAY"	S	g�) �V��@ ���	C&� 4�  ���T	�j�H���J���3�]��@-�S�Qb� g� bN�2RT
�
�p�����%? ���$?�%-'>� B�#�E�Y�0-5�S��s�3�h���x� (�'&�>�U`�t�4��^�R`�	U
 	pZ���� ��@dr�&�E��@<�E1su�KP��U���ԃ>c$B���@����	��%v2Ӏ��% ���;�tȠ�����-�e��	��*ȴ��F� (��f
�u� b�� ~]v��U�m��8S�	)��*[r����_�r���+�'�: ��'�!J�ԢLu���.�y��V,�Tl�w/Cf����$��w����wHT��T ݠ��<�s<����o*��A �>�Ct�F ��&�� ���t�&���&��w�+�:�P=Ɗ $<@w�:�9v�2<�<?w�+����)�,$H�! �<�3^�I�f�@� �4� @B�, B��P���Èw�%HID�]�G(����%�����������3ۇf�tX1�>�!xsHCPrXaM�0��u;M�A�PA��5	��-:P��u'��x\W<! *cD�_aT�����bR"!	xucY4U
a)Rt�J!g:)`ta('ģ�|�4����Ĉ�bn4oe�u�,"�"E�� �ب	= s�K�+}�F�	����MV�T,U�?�bA����Ro���LJ�Ɩ$eJ�$�$$tI�$a$E��
�@�LZY�	��"-:  SR�>0 u/3�K�� 8�A��2�!
U�6
J��4.t�5*� #Z��<O�O*@8�v��\�T ��u�X�.Rt\�\iH��.�%PR���  bZX.�>��t1�<t P�<
t�<t<u�
$.(s�.�0 
 P�1���u�u��X�C23�S06� �[ͥ3&L�T�F�.�.� G	�PV��.�Fc<�p����^1��e�P��
�`�E=�0�<t��/I�����3��� �5����
�<��t= rt��Vl�u�5���.����6,�Ŋ���6Eb�Hs7�\�R�(��^�Zcw2��1`\� \�
����  �{�r���=t:��t �< |��s� C��B*u	Q4QEQ�k� �K����z
�
u�����8�* z���) 
�[+��`d ^c
n 0GETLINE BUFFE�@  �8<zw, �9�� }uF��Æ�� �  �� �Q�PX��P$  <	v0����u�X Y@RWU����5�0� �h.
z��%O�`��v�G����Y��]=_Z[ڹ �';�r���������1��� �
 �DW��0�X�����P�P����=?�=�d �{�����d���=��
�xV��6 ��8@tV$�4��^Z�Q$Q�F:�t�C��1F�ܷ P���0r'q	w"� 1�<<bt(<w  t*<at,<tt2<dt=<r t?<ltFP�@���X �9����륓����Rd���R�����R�C�@P;�Z��)���#�
 ��R�Ĵ ,0��D��������%�P�W� P@$���H�r!��K>�$ � ��3������V�������mRV5\*����X00 @t���r�D<Dt�T�����F��� ru���#
���H �ʀ� ����^�z%z��d����K��q�;�v"� Q���� ��V�")�>*�L)��^������q��L���@���t*�(�<2�(�0��������ݝ)���������Q�>4�2xt=� �2FC � ���`��0�F
V�4/G �.7MSG 
=)!.i�/0	��
& [�%�q�@<a� �nF�	��P  *rr-%�5Wб@� �6�		�������a ���
<r�pt ,� �5��L�ffH�}��� �#�m��à �s��H��Þ���p�t9����v�K������O�&� �M�&��0V���R�S� � rK</u�N�}� A��?��~�G�u������8	�����R ���+�v!�����(� B|�������g� �.��O� �	@j��:�}����_����(�(f���G�� �~vP�<,t	�� �S���&Y��!V�ߍ7IE4I�b�� X@}t����w�o�.��l��E�V (
Are yo��u su	wantP�*o dthis?((#Ifo, p!�$ss Y; !ynPJg els4cc*�	.(? N|YTJ0nrDd�=kI7buiT�ld 2riv��2@0a:&7d�0SENTuT!whe!ady�
K�   JCAUTION !!T��{ttempts�XcoNrlY�l�Wfe�0N los{aftB5form���gum))��'�no%�9bequs��?�T�Tm2�.)�qmeod�@3guarMU9'po/L
�y of]�r��AR�s�rch-pha@*+Ps���e:A�1�l��Non��@5=Y��@Il�%V!l%#agaP�D�UY�RA��@_wri�AoDD�,Inv`i]�(�unsp�i�vI�. ɂ�r��DOS ��s�t�C�{c��n�w��)k9Yp1(s)ѫFAT�8b�O'd�RoL�i�{Fy$=A�plac<P3#Simu�@�Fly	�a�, #ST,���gnizR4 N6e! ;ugh�mϲrBc�a`take!�� sys��a_�KEr~([f@1&s�#U2w@3wh~Bwd4@�5t+G� �d�e-�U�;bf*��#  ΋vyEկda��<s$qu!Eeru��C�E��ek
Lk"�Hwn�wa {��[f�Y1N���pO���aul��F�gen alLvil_^ �"f�  <��>F
VO!L
ExaҀi@0�oB�f�i��%�{�z%�4�":x,�ub�� i(S%CmY�.�K[%
��~, 1���OyM.�:*@�_1d,{��Uzm5
#�mr�.�,�* C(6R�bxulx� *Walk�+� �t	C e�loca0��P�Y.PC��.c7k,ragm,9U	�A'DpeP
% c�ssl
k�~-O�!+�\zNytH)��ab"��!Tr�}bm�Jef�A? ��!�SH�sM���9H�rn�!  � nex�e}pXs:��q�8
��6sg	�]O���]�E
Ewsh/m5dn9��� (YJH/No/Qu�)"��Ign�0���q� KP��ut{:F!L&PT1gR$li���h�t`�s� B�FORM/ݪ�GN+~@�&RECOVER5/N ��eUN=@'y: [/J]
U]ͱLO��P(��#��V 9S�s\!�9��un9.��-�[� V�,��1mi�ag���wie�iK���M���fup U�1sKG�y����:_2�|3 LD.�@# e< Inam�M�,�hu�~���A
,sc�p��iAy�u�)���b�N��N D/� b���do�kaP���z�SZhd\2�6p9�sa+p����cUn��ƿ ��>.�v�	�

(L�UNDELE�,5�(0Copykgh~ E(C) 1987-93�#�Po��ofB�tw7,dI�c+i�h=@0t\U�%���@ H-d"�͔P�T�%o���ph�?,>rw��[B:
t[�@l� \�agtype�:  ttq��C�W�p? A�+��O�^"�6mp���s: .{#.����^ε�H:f��Ҋ;x�z,=$$r70D}/d!Pxװ RsW�S���=�-i/��" �RU�?R�\ �2)|i`�`2;�deX�kippf7�v t��vwasa��D��7�a��l�i6�-��#@�(DL=�bh):��J,�Q=�Y�,i���#Y�.�1/Y(Bhw� ��s��{9-�?��;�=l� ��H.�A�~A�8�Whi~ԉ�?� **�e (BQ�I�,q1�8CylB����Ԋ�3-|RbU{a+G�b�f���A ���F��&����d��K�0�`����+d��r�3d�r&(4�Nt���" [�f�dollowǏ8q�oF1�4b�P���r,dm,�tn:u]�Ta��al_�˪�4��_ �E��X BT�ӑBJ�~�T��C̳� H�R$l#z�M- -����OS16 2`HUGE���XTEND B� �� RP? oUJra�;)l��6r)l��4<���`�signa�|��]���Z~q`v��C�p�im!��c*֕�GZV� �WARNINGÃX�~� �'�#��s�i����6�acq�J��d4bt&f�*�I�� �"��n�tEr�'>'|Y� s'ca#����h#y��;}mod逆#ce	�+�,]�w09�U�=��%��J}B�2$$`auhb '�(_w�X�m!Neq��p 2.x��og�#�b$c�{������iBa���bypa�� T��6&�t�Z�n2P�s���.Z. It/��R���ic�Eb��bat�lt$F*	�vJC$ vm�6�59���P	�XX:� DMM/DD�m/YY]f6�up�� Tp(Y/ѠN$
JOn��eGF��zr����x���7���_ñk� �nGe�ٕaΆ�H 9�Xv�٢ IjC���JW�o<?	�90@Ifi�miWsj\u��kdic�Ԙ+��
LL��k?K��A �@P@P�}pSC󬟌^b5�ny��O(��8�oZ�7 �x�3��-ˤ�
�ry�)RDkEs%���1��mN 7m ������ =zlog�l�_� s�,	 A=AЂ�xR=ReR��y	I=�!�e!c%hO��U w�Ra9� x }a��W7GY"D�.Z�Inuy�UO� t,a3�ckup�mo8��D1q�
DM�o�sqᖭ鷼�o��-�gˋ���7YBĬ�ke�O�3�� X� �E�BAKV�
��9x:\��5aMS��ESLIFVASIM0�AEP��
REB�8UBD`$0@.$.��<A.��<Q��6M8�
9.���  =A�� �� t.�-=(
��W!��	� �!�S$0=s�� �+u|�\l`rJ8 � r���@ra�e�>.= w۝�83�x�� `�R.��(�k7C>
u��464uM� <7<�{6Dv1>P�4�X��9t�ws�s.�#=.���|��%~<�r�
�.�8�.j�~TI*Y>�6 ��� �0�R@/�;n<t"�� u�<R����e�� �B�p<u��J�r��J�t��J%v�k9E��u����u��(�����<;�%�"���{v'�@p��<;�v���V��&���.0>�s�O.ŹuJ��E�E:4+Ecr p��ìt�w;p3����9Q �<t$�< XLt<Pt����DY7��(��2ӝ7�7R;ut)8G0GN~��Yu� :�@ �\�Rl.��r��ܑ<����,dk7���,�G(s �&�v(r�3��Fp:u�G,��++��.n8>8�(����NQG�hC�.J� ؂V���M J6k�.��<tD."�+.����������G$�r!:@Mu���33W������>=�u	��d� �X��7�R��I���=-l#)��38S�!2&[28�{ 8D��7�Ńm �j'r:8�j'9u8�j)jN��j+2���j+2��zjj�j�b�4.����/2 d�8= w3.�6N�EK<����bY����PS�g�or�?b�2!4Ǖ  (�F)����|(�[X���ø3�
 :���r���� 0��=u��u��b1=�T@t\��L.�x-z�z�� 7@����Tɣ`����T�l�=�S��� ��rR�
r�,.��$*  $9	s%){0�>vn�a tBh� j�6 KcK ,�s�R���eRZ�Jir)�&�6k9*9���gr����	2�$�u�x\�<u8B�":�!�
�Yt<Nu�O���s��[�x)/�z<~�	��� s8�
 ���Xy.�Wy�<r����B�]� CU3� =Y5(I=�C_;I)EaG�c�I�e;�Pp2;��>�� �������;�ҋ�����U�˼+�`(��S-:� l<��.�<�� ��e��[�(�>��  X�uFGI�uz�u�P��,���ދDك��<=� 1j�� D.�T
!(|! uRrB|�i
�M�9D!r		|ā	w)�
J2�#9%�!%''TR#)%1+=�V 
p�< �2.����@���� ! �r�>1= ��� �x�trPRS�D11�1[r
<uh�O.��	x�@
� +Htj��u�C��r<�pT��P��* 	 =XH� �O(A��(g�g��n<�G��@)5��@ZlI�v<��.�!�.�&�f��t������6�� ��^�0�SQRVWU�#��������I.�y5=
ꋠ�,�DA�Rt�`��5 �%r
��]_^ZY,[Ýu�� a�  � r��I1��"��C;u&ut��u�F��:=��������0�C=h"   At<Rt
<IuY��XO3�8 N>��� P$X���0WVQP.�>���6>n� �t��% =	�
�9��+�� s� '.=XY^_�VW�Q�� ��A�V���^(t=�<v��( �Y��RS3һ
  ����00[Z@�YQRWU��3� CH�bOC�EG�>I=�'8���C�Em�q��K� ��0�O�u� t���#�3�3��h�]_IX�
�7P"�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              ���ó\-+|                                                                                                                                                                                                                                        \                                                                                                                                                                                                                                                                         
*.*               :.                                                                                                                                             ������ �����Ns
����@���!��A��� �6 �F r �����A�´G�!�@�� ��u��������L�!� � ���r�>�������	� ��	  �r+�> u	������ r�> u��\���� �G�!�Ê:�t(�
�u��A��!��!:��u�� ������ú}��!� ��/
�t���/=��u����/��$5�!�y�{�*	�$%�!�#5�!�u�w���#%�!��3��/�P���}����,@��QS�?� � ���C��[Y�}��!
�Xt	�������F��� 󤿩�m� ��? �5��� �,� ��N�!÷ ���@�� i�!r���������&�PW������ �+���I_X�U��o���-!= rl�>\t(��;�!r���@�v.�F-\�G�!�v-��A ����~-�A ��;�!r�A��t�E ��g�� ���������� �����o]���u��F+���F+À&��������!�  ��N�!r������<�O�!s��r�� ��� �$����!�rc��$tP�>�.tI���}��� ��L ������ �+ ��F,������� ���+ �F,��.�V-�;�!�>� u�~ 뛀>� u�þ� �G�!N� ����\t�\G��� ��3Ҭ< t�1sF� �����Nú���!� ��N�!��O�!r�&�����r��$t�>�.t�����u1���}�+ �O�!r�&�����r��$t�>�.t�������� .tD���@ �k �~ �/����t� � �F+�>��.���$t� �>��/� � �Ë>��$u��2���2� ��� ��< t��O�
�2��Ê�$u�+ �F+�>��.�Ê�$u� � ��� �>��/�à8F+u�F+ ��8F+u��F+�� u���- �S� �@�![�� = u������SQ�  �Y�!Y[�SQRV��]�u�M�U�s���]�u�M�U��^ZY[�� �L�!� �u�@t���;�!����!�t	����/�u�#%�!�y�$%�!�P�.�y<|X�&��A:�u����L�!���V�6�uP� c�!&�6&�X�< t:r:Dw�������^�         �	  �	�	�	  �	�	  �         �	�	/F /A �          �	�	/?         ���	=  t� ���6�	� r�>�	�6�	3ҋ�	�=��u��Ëځ��	uL�6�	�|:u
�>��FG��>V���^�@ A���< u��\u��\t
��@ t�E� ��
��>��L���4�>�	�	u�N ��&��	=�	u��	 �����	 ���	�ã���	;�t� ������� �>����Í>����>/t����                                                                                                                                                                    �    �    []|<>+=;" ��
  ���
��
  ��
  ��
  ��[]��|<��>+��=;�s���S&�&:s� [��6�
SWU��
��
 u>��#r7�t2�u��
 u�W�"��
AtN��<=u��
C�sɬ�C��N�6�
� ��
&��6�
�</t1�<"t��
uP&�G2�9�
s��
��CC�&�� �f��
 �^&�G2�@���&�2��tCS&�� [s?CC����
 �3&�G2�@���&�2���@�&�2��tCS&��T [s
CC����
 ]_[��
��
�6�
��
��
��P&�� u��
�< u� u��
 �P���� X��X���UQ&�O2��t�o	�s� �����.�
�Y]�&�~  tE��EÀ�
���rB�&�
�P��
+��
X�6�
�< u#�|�:u��
	 �&�? t&� u��
 �	� ����
P���� X��W&��>�
&�&�eP��
&�EX<u
&�U&�M�Y<u&�U�O<t�<t�<u&�U�=<u��
@&�E&�]�+&�u&�]P&�Gt��	&�Gt�� X&�Gt�d _��� P&��uPSRW��
	 ����`�_Z[X���$�� t��
  ��>�
	u�  t	��
  � �>�u�>�
 u��
	 X�PV�
�t<:u�| u� �	�sFF��^X�VR�Њ�}r
�t� ��FF��Z^�<�s<arB<zw>$��:SW�>|��t�>w8tPQR�e�»��� ����!ZYX�]�ECC,�&�_[�<0r<9w,0����PSRW&�&�
�u�����
	 ����c�_Z[X�PURV����r:�r���
t<=u&�~ un���
t<:u
&�~  uZF�Z&:F u
�tPFE�&:F uCF�E&:F u9FE���
@t&�G  t&�~  t"&� t<:u	&�~  u�< u&�~ :t���6�
�^Z]X�PWV�>�
�
�t�W u ��^� _�9^� _&� u-��
 �%XV�
�t�* t�sGFGF���
� G�>�
^_X� t	P����\�X�SQ���	 :tC��AY[ì�  t�Q u��
 t���
At	N����N���SQ<t-< t)<
t%&�}r3�&�]��&�9 t3�&�	C&:t��<Y[�SQ��
 �&�
�< t6<	t2<,t1< u�< u� F:��&�}r3�&�M�t� C&:t��< Y[â�
��
u��
 :���.�
;�t
</u����
</u��
@��VS�>�
 u%PQRWU3��޸ c�!���]_ZYXt%�6�
��
�6�
��
�< t:r:Dw��FF���[^�                        �          �  � �           �       �  �  �        �  �     �0     �0,      �� ,  @  c  x  �  �  � ,� -� ./OIncorrect DOS version
&Directory PATH listing for Volume %1
Directory PATH listing
No sub-directories exist

Invalid path
Volume Serial Number is %1-%2
��óDGraphically displays the directory structure of a drive or path.

!TREE [drive:][path] [/F] [/A]

;  /F   Displays the names of the files in each directory.
3  /A   Uses ASCII instead of extended characters.
�>������ Extended Error %1�>��� ��� Parse Error %1�>����            ����        ����        ��������    ����       
     
 $$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$MS DOS Version 6 (C)Copyright 1981-1994 Microsoft Corp Licensed Material - Property of Microsoft All rights reserved PSRW3Ɏ�3��.� �/��>�.��/�"�> �.��/�2�>0�.��/��>����>�.�>,���&�>$�.��/�:�>8�K
��$�P  �R
 �(��><� �. �A Q�P rY_Z[X�����PV� c�!r�6D�F^Xø D�  3��!�����D�!ø D� 3��!���D�!ô0�!=u��= s����� � �  � ����PWU� r����t���]_X�VS3�3ɀ��u��<���%��tļ ���= r=' wļ,���ļ�Ã��u���u���P���� 3����� t�T ���r�u럜��u)RUQWP� �/<�Xu	�ظ�/��s_Y���� ]Z�����[^�WP���2����IX_Ã�u�>8�t=��uP�P�8X��8�3ɀ��t&�M�	.85u.�M���s-��t���t&;�.;u�	It�����r����u&}r2�&�G�J �PSQUWR��H�6M����t�u�& ��rZ�_�����_Z�r]Y[X�����PSR�H���u�, ��w s�Y�  �!2�������t;�t� ���rZ[X���u�&��!��� s&�U�!����t	&��!GIu���WPS���ٰ��u+�K��[X_�3��tO�@�׃�u(�!P&��Z Xs��@B�!�&�=u��������UQ����Y�!s�;�t;��u��]ø' � �À��t�ƀu�>K� � ��W�>D�t&�= �t&:r&:Ew�GG��_ÏN3ۓ��6R��6R��	v��7���0RA�u�t9��u�|
,u�6[A�"��u�|
,u�6[A���u�|
,u�6[A�3��3�3��6N�3��t!�%� &8%u
&8et:�u&��S�sGGBIu�V���t3M�>P u+�D0&:Eu�<0u�t4��>M�uBBIIOO����W+��
�_Ys��Q�ʀ| t�tIIGG�^��u^�	���u3��tVUWQ3Ƀ>P u-�Du�|�L��Dt�Dt�Du�|�Z� �R ��  rY_]^���
��>P ur���P  �3ҡP�R
 ��X��TC��@u�� ��u�
��TCC�� �3ۀ| uǇT -CCƇT C� ]3�3҈J�D	:�v*����D�t�D
��TC��@u�| ��u�| t8Ls*L�ъL�t$�Du�Dt&�G�X��TC��@u�A ��u��D�u
�t�D
��TC��@u�# ��u��Du�Dt�
�t�N��u�� U�QW��3ۍ>T��r_Y�����]�D0u&�PA�h�s&�EP��&�
�tGA��+�U�]3�3��R 3��D u$&��Du��tC$�R
 �Du�R
 �T�Du&&��Du�ĀtC���R
 �Du�R
 �(&�&�U�Du�ƀtC���R
 �Du�R
 �D@t)PR�82��T�!s�[,�D
��ZX�D
,����ǈD
�����t3Ҳ-RU�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               MZr      M����    r                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      � � ��    �    []|<>+=;" .�   �.� .�   .�   .�	   .�� [].�� |<.�� >+.�� =;�os���S&�&:s� [�#.�6 SWU� .�  uC���r<�ct7�u.�  u�+�&.� AtN�.�<=u.� C��sŬ.�C�N.�6 .� .� &��6 .�</t6.�<"t.� uT&�G2�.9 s.� ��CC�&�� �i.�  �`&�G2�@���&�2��tCS&��� [sACC��.�  �4&�G2�@���&�2���@�&�2��tCS&��] [sCC��.�  ]_[.� .� .�6 .�	 .� ��P&�� u.� .�< u� u	.�  �P���� X��X���UQ&�O2��t�o	�Os� ����.�. �Y]�&�~  tE��E�.� ���rJ.�& �P.� +�. X.�6 .�< u&.�|�:u	.� 	 �&�? t&� u.�  �	� ����
P���� X��W&�.�>	 &�&�eP.� &�EX<u
&�U&�M�Z<u&�U�P<t�<t�<u&�U�><u.� @&�E&�]�+&�u&�MP&�Gt��	&�Gt�� X&�Gt� _�.��  P&��uPSRW.� 	 ����[�_Z[X���>�� t.�   �(.�> 	u&�� t.�   �.�> 	u�  t
.�   � .�>� u.�>  u.� 	 X�PV.�
�t<:u.�| u.� �	�%sFF��^X�VR��.��r
�t� .��FF��Z^�<�s<arE<zwA$��=SW�>� ��t�>� .8tPQR�e�»��� ����!ZYX.�].�ECC,�&�_[�<0r<9w,0����PSRW&�&�
�u���	.� 	 ����8�_Z[X�PURV�.��or<�m�.� t<=u&�~ uq�.� t<:u
&�~  u\F�\&:F u
�tRFE�&:F uEF.�E&:F u:FE�.� @t&�G  t&�~  t"&� t<:u	&�~  u�< u&�~ :t��.�6 �^Z]X�PSV.� �<"u!C�/ r.�D ��F�� .�6 �.�6 .� .� 	 ���	^[�Q�X�P��� t$<"u��"u.�FCC���{s.�FC�.�FC����.� �X�PWV.�> .�
�t�_ u$.�� ^.� _�?^.� _&� u2.�  �)XV.�
�t�- t�sGFGF��.� .� G.�> ^_X� t	P�����X�SQ�� �	 .:tC��AY[ì�" t�S u.�  t�.� At	N����N���SQ<t-< t)<
t%&�}r3�&�]��&�9 t3�&�	C&:t��<Y[�SQ.�  .�& �< t6<	t2<,t1< u�< u� F:��&�}r3�&�M�t� C&:t��< Y[�.� .� u.�  :���. ;�t
</u����</u.� @��VS.�>  u'PQRWU3��޸ c�!���]_ZYXt).�6 .� .�6 .� �< t:r:Dw��FF���[^���  �: [ �  � �  ����� �  ����� �  �� �    ����       
     
  �$A �MS DOS Version 6 (C)Copyright 1981-1994 Microsoft Corp Licensed Material - Property of Microsoft All rights reserved v � 	 �  �;�;���   ���  �   		  		    		/N /V /C /I /?K �  �
� 8  L  ^ ,a -� .� /0U1�2�345L6�Incorrect DOS version
Insufficient memory
FIND: 2Searches for a text string in a file or files.

DFIND [/V] [/C] [/N] [/I] "string" [[drive:][path]filename[ ...]]

E  /V� �  �Displays all lines NOT containing the specified string.
E  /C> �  �Displays only the count of lines containing the string.
=  /N> �  �Displays line numbers with the displayed lines.
K  /I6 �  �Ignores the case of characters when searching for the string.
0  "string"  Specifies the text string to find.
  [drive:][path]filename
4� �  �Specifies a file or files to search.

LIf a pathname is not specified, FIND searches the text typed at the prompt
 or piped from another command.
�>	������ Extended Error %1�>�� ��� Parse Error %1�>1���PSRW3Ɏ�3��.� �/.��.�>��.��/.��.�>��.��/.��.�>��.��/.��.�>���.��.�>�.��.�>���.��.�>��.��/.��.�>�.��
.�7$.��  .��
 ��.�>�� �- Q�< rY_Z[X�����PV� c�!r
.�6�.��^Xø D� 3��!���D�!ô0�!=u��= s����� � �  � ����PSQUWR��.��.�6����t�u�& ��rZ�_�����_Z�r]Y[X�����PSR.�����u�, ��w s�Y�  �!2�������t;�t� ���rZ[X���u�&��!��� s&�U�!����t	&��!GIu���WPS���ٰ��u+�K��[X_�3��tO�@�׃�u(�!P&��Z Xs��@B�!�&�=u��������UQ����Y�!s�;�t;��u��]ø' � �À��t�ƀu�>�� ����W.�>��t&�= �t&:r&:Ew�GG��_�.��3ۓ�.�6��.�6���	v��7���0RA�u�t<��u�|
,u.�6�A�$��u�|
,u.�6�A���u�|
,u.�6�A�3��3�3�.�6��3��t!�%� &8%u
&8et:�u&��K�sGGBIu�V���t5M.�>� u,�D0&:Eu�<0u�t4��.�>��uBBIIOO����W+����_Ys�g�Q�ʀ| t�tIIGG�^��u^�	���u3��t>UWQ3�.�>� u�Du�|�q� ���" rY_]^���
�.�>� ur�*�.��  �3�.��.��
 ��X.���C��@u�
��u�
.���CC���VS3�3ɀ��u	.������(��t	.ļ����= r=' w	.ļ����.ļ��Ã��u���u��.������ 3����� t�T ���r�u뚜��u)RUQWP� �/<�Xu	�ظ�/��s_Y���� ]Z�����[^�WP���2����IX_Ã�u!.�>��t=��uP.��.��X�.���3ɀ��t&�M�	.85u.�M���s-��t���t&;�.;u�	It�����r����u&}r2�&�G.�� �3ۀ| u.Ǉ� -CC.Ƈ� C� ]3�3�.���D	:�v*����D�t�D
.���C��@u� ��u�| t8Ls*L�ъL�t%�Du�Dt&�G�X.���C��@u�C ��u��D�u
�t�D
.���C��@u�$ ��u��Du�Dt�
�t	.����u�� U�QW��3ۍ>��Q�r_Y�����]�D0u&�PA�8�s&�EP��&�
�tGA��+�UÌȎ�����s��������=�b�!�۾� 3�.�	�>�  u� �� .�	 �O&�	�!&��t�9�7&�	�~V�	�>�3�������t-�e���� �����!G�=&�� +ã����>����>	�t3�����=� �!r]P�>	 t'��(��(2��
��������u	�	� ��X�غ�� �?�!s�;�u��t�#�u�w�>�!�]�)WQ���Ȍ؎����uO��+�Y_�t�S��P�Ȱ
���X��u=��݀y�
t�G�
GWU��J�� ]��Y�ٰ
���u�QW��+͋�I&�}�uI���a��RZRB�W����_s���v+;t*��:t$��t	�%�A:�tXP@+�+���nr��Z�JJt�`r���� Z��t�z���u�p���t���b�R��t� �Ջ�� Z�L���[�t�ڹ����B�!r��#�tM�>�!� �= u� �� ����������� � ��]��^.�	�.�>	�t����9.�� .�� �S#�t	��� �3 �����2 ���$ �	� � [�SR����� �]AA��� Z[û �@�!û
 3�A;�r
3����0R��0P��X������<�r�  ��<�r� <ar<zw$߆�<ar<zw$��SW�>���2�+�&�_[���S sGI�GI����WPSQR�Ȏ����e����� ����!G&�.����&�.������&�.��.��ZY[X_�VP�6������&�< u��&:s�&:Dv�����X^ôL.���!���� ���ÿ�3��4�=��u.�	�.�>	�u_��#�t��1.�>		t%.�>	u.�>	.�	��7.�>	t��
 ��.�>	�u�
 ��� .�>	��� .��.�	��.�>	�t� ���� �PSQRWV��3���=��u� = u� �� #�u�.�>		t�.�>	t�.�>	u�.�	���u.��봁��u.��릁��u.��똁��u.��늁� 	u.���,� 3ɶ����=6t@���� ��# ^_ZY[X�.�>	�tPR��� 3ɻ ��ZX����3�.��� �����WSR3�&��t&�C"�t<tBG��Z[_Ó� ��
 �-
 �  � ��������    R���RB��� �  ��� ��O����P�4 PˌÌ�H�؎�� � ���G����H��� ��������+�s��+�����ڋ������+�s��+�����¬��N���F��$�<�u���<�um�¨t��2� �3ҭ�����Î�������t&��� �t�� �܌�@����&H����Ë> �6
 � - �؎��  ��֋����.�/�@� � �ʎں�!��L�!Packed file is corrupt                                M�DOEQ$ESDEUdEW�EY�E[�E]�E_Fa$FcDFedFg�Fi�Fk�Fm�FoGq$GsDGudGw�Gy�G{�G}�GH�$H�DH�dH��H��H��H��H�I�$I�DI�dI��I��I��I��I�J�$J�DJ�dJ��J��J��J��J�K�$K�DK�dK��K��K��K��K�L�$L�DL�dLǄLɤL��L��L�M�$M�DM�dMׄM٤M�����M�N�$N�DN�dN�N�N��N��N�O�$O�DO�dO��O��O��O��O����/PEPeP�P	�P�P�PQ%QEQeQ�Q�Q�Q�QR!%R#ER%eR'�R)�R+�R-�R/S1%S3ES5eS7�S9�������S?TA%TCETEeTG�TI�TK�TM�TOUQ%USEUUe                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                MZ�K     ���	�    	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      U��$ �-j�F�P�F�P��e���F�t�F�P�F�P�/f����P����v�v� �����  RP�F�P�F�P� P� P�6�F���  RP�F�P�F�P� P� P�6�F���6�R"P��P�  P��P��P��*�P�`P����� P� P�� P����= u �� P+�PP� P� P����
� P�i��+�P�`��]�U�츠 �;iWV�F��v�v����Ɔ`� �F� �/�^���v�0��`�P��|���F9F�t�� P��`�P��|���F��F9F�~ɸ� P��`�P�|���FH= } �� P+�PP� P� P�4��
�W P����FH= } �� P+�PP� P� P���
�W P����^�_��P��d���^�_�Ȋ�P����d��;�uA�^�_�:u5�^�_� u)�^�_�:u�� P+�PP� PP���
�W P�$�����`��F��F�  � �F�  �F�* �F�P�F�P�!R���F�  ��^��v����<	�F��F��F�9F�r�^�Ƈ<	 �~��v�� �~� t�~��u�F� ��F� � P�v�� ���~� t!�9F�t��9F�t�9F�u	�v������ �~� t�[��^�w��{��= r	�v�2���v����v�v����^_��]�U��3��(gV��^�7�</u�|?u	�| u�v �N�F�~ u�^]�U��3���f�<	��� �� P�J{�����~t�~u�F*�P+�P��F*�P+�P� P� P�v���
�W P���]�U�� �f�F�,�� P+�PP� P�v�����
�F��~�:~�+�P�h��]�U��3��Wf�~3w�~�s�� P� P�B����~w�~s�� P� P�(����~w�~s�� P� P�����~v&�~t�~t�~	t�~u�� P� P������~u.�~v�� P� P������Ft�~v�� P� P����]�U��3��e�~v�� P� P�����~<r�� P� P�|����~<r�� P� P�h���]�3��Ze�* z�, �- �. ;�/  �z�{�|�	�~�	����������������  ��	 ��	  ��	�	��	�	��	 ��	  ��	  ��	�	��	�	��	 �� ��  ������	���� P��P�x���� P��P�x���� P��P�x���� ��  �����	���� P��P�nx���� P��P�`x���� P��P�Rx����  ��  �����	���� P��P�'x���� P��P�x���� P��P�x���� P��P��w���� P��P��w����  ��  �����	���� P��P��w���R"  �T"  �V"  �^"  �`"  �b"  �X"  �Z"  �\"  �d"  �f"  �h"  �j"  �l"  �n"  �p"  �r"  �t"  ������� � � � �U�츐 �c�F�!e�^�G�F��w��p�P�
w����p�P�]w���F��F�P�F�P�x���^�w��p�P��v����p��F���� PS��v���u�� �� P�v���v���u� �P�v���v���u� �P�v��v���u� �P�v��v���tw�P�v��v���tf�P�v��v���tU�P�v��wv���tD� P�v��fv���t3�%P�v��Uv���t"�*P�v��Dv���t�/P�v��3v���uD�F��� �� P�@v����� P+�P� P� P�
 P�,��
�W P����F��^��? t�����]�U��0 �a�F� �^�_��P��]���^�_��^�_��F�<A|<Z�^�_�:u�^�_� t �� P+�PP� P� P���
� P�+���^�_��`�� �� :��  �� P�F�P�F�P+�PPP� P�P+�PP�!6�F��t �� P+�PP� P� P�E��
� P�����~��v�F��؉F��N��F�D�F��F�F؍F�P�F�P��u���~� t@�F�D�F�	�F�F؍F�P�F�P�u���~� t�F։F��!�F�  �F�% = �A�N���FֈF��F�  �~� t �� P+�PP� P� P���
� P�#���~� t+�P� P�� P�e��� �F�+ҹ
 ��0�F�F�+����0�V��F� �`�F��F� �F��� ��F�P�/t�����F�	���F�P�t������ P+�P� PP� P����
�� P� P+�P� P�
 P����
�F�D�� ,@�F�F�P�F�P�t����]�U����B_Vǆ�A ǆh� �F�!e�^�G�F��w�F�P�-s���F�P�s���F�F�P�F�P�8t���^�_�:u�^�_����<A|<Z~��x�P��Z�P��6��x�@����^�_����^�G���B �C :�D  8`u�� P+�PP� PP���
�W P����B P����P���P+�PPP� P�P+�PP�!6�F��t �� P+�PP� P� P���
� P�8�������v�����؉�������Ɔk�DƆj�������l���j�P��j�P�2s����v� tIƆk�DƆj�	������l���j�P��j�P�	s����v� t	��j��F��#�F�  ��p�% = �A�N����j��F��F�  �~� t �� P+�PP� P� P����
� P����~� u[���F��F� �F��� ��F�P�q������ P+�P� P� P�	 P���
�� P� P+�P� P�
 P���
�F�D�B ,@�F��F�P�F�P�4r����*�-@ �F�P��^�P���P�;6�F��t �� P+�PP� P� P�=��
� P�����^�P�q��= t/�4P���P�p����^�P���P�[p�����P��^�P�p���^�_�:u=�^�_����<A|-<Z)�~t#� P+�PP� P�
 P���
�W P�:����^�_����</t

�t�~u��^�P���P�p���6P�� ǆ�  �����^�_���� ���</t
�u�^�w���</u� Ɔf� �^�_�?\u�^�_�\t�^�_�?:u � P+�PP� P�
 P���
�W P�
���^�_�?\u�^�w���P�xo�=��^�P���P�io����^�P�o��= t�;P���P�
o���^�w���P��n�����P�o�����ǆ�  ����������.t��� uꋶ����.u���.u���\t��� u�F� �������9��r�����������������\u��P�F�P�n������B� ǆ�  ��������z�*t�z� u싶��z�*u#�� P+�P� P� P� P��
��
�W P�T	���~� t�N����z�Ɔ{�:Ɔ|� ��� u�=��F�P��z�P��m����z�P�Rp���tD�^�G��� ��w�^n������ P+�P� P� P� P�J
��
�W P����ǆ�A �vꍆ��P���P�;6�F��tP�b
���v���������Ɔ�:Ɔ� ��^�P���P�Em�����P�o������P��m��= t/�?P���P�[m������P���P�m�����P����P�;m���AP����P��l��������P����P��l������P���P�m�����P�[m����������\u�CP���P�l����f� u�^�_���� /�^���G�����Ɔ�:Ɔ� ��^�P���P�bl�����P�B P�l����P�  P��P��P���P���
��P��l��= v��  P�l��= v�� ��P�l��=@ v�� �GP��P�fl���u�� �LP��P�Ql���u� �QP��P�<l���u� �UP��P�'l���u� �YP��P�l���t~�]P��P� l���tl�aP��P��k���tZ�gP��P��k���tH�mP��P��k���t6�rP��P�k���t$�wP��P�k���t�|P��P�k���uD����� �� P�k����� P+�P� P� P�
 P���
�W P����F��$���*t���?u+�P� P�� P�B����F�^����
�u�^��]�U��3���V�9Ft�� ��;u���;u+�P� P�� P������;u"+�P� P�� P����+�P�  P�� P������;u"+�P�@ P�� P���+�P�  P�� P�����;u"+�P�� P�� P���+�P�  P�� P�q����;u+�P� P�� P�W���9Ft�� �*�P�P�P�5�����;u6�*�R"��T"��V"+�P� P�� P�
��+�P�  P�� P������;u6�*�^"��`"��b"+�P�  P�� P����+�P�  P�� P�����;u6�*�X"��Z"��\"+�P� P�� P���+�P�  P�� P�{����9Ft�� ��*�P��P�6������;�u6���d"��*�f"���h"+�P� P�� P�.��+�P�  P�� P�����;�u6���j"��*�l"���n"+�P� P�� P�� ��+�P�  P�� P�� ����;�u6���p"��*�r"���t"+�P� P�� P� ��+�P�  P�� P� ��]�U�� �3T�F� ��F�P�F�P�/ P��h���~� u��  �)�F���F�P�F�P�/ P�h���~��u�� ��� �>� u9�F���F�P�F�P�/ P�h���F���	�F���F�  �F�P�F�P�/ P�ah����]�U�� �S�F�t= t= t"��P�s���%�^�F��^�F�� ��^�"F�F�
�u� �+���]�U�� �CSV�v�g���F���N��\ P�v��v����u�/ P�v��v�����tՋF�F�F��F9F�u�؊�F�<\t</t�� �^�� �v�v��f���F�  ��v�v�</u�\�F��v�$g��;F�w�^�? u��PS�f���^��\�F��v��v�f���^�?.u)� u#��P�v�~f����P�v
�qf����P�v�>�F��F���F��^���F�<.t
�u�?.u&� �v��v�9f���^��.�F��v��v
�$f����v�v�f���^
� ^��]�U�� ��Q�F�����~� v�n� �v��F�P+�P�K6�F��u݃~� t'�~� w �� P+�PP� P� P���
� P� ���F��^�\  �~� u	�^�����^�F���G  ��]�U�� �cQ�F� � P��P+�P�K6�F��t �� P+�PP� P� P���
� P�. �����f�d  �^�F����]�U��3��Q�v� ��]�U��3���P�v�����]�U�� ��P�B P�g���� P�g���~ u� P�@ P�� P�����u�F  �F�t= t=  t=t��F  ��F ��F ��F ��F �>� u�F����	�F�F�P�F�P�/ P�e���v�uO��]�U�� �:P+��F��F�� P�� P�� P�����t� �6��6��	P�v��v���6�F��tQ��	P+�P�v��v���6�F��tP� ���v��������	P�v��v���6�F��tP�w ���v������� P+�PP� P� P� ��
�P����]�U�� �~O�F�F�F�F�F�F��F�F��F
�F��u*�F����F��F�P�F�P�hK�F�u��]�U��3��5O�� P+�PP� P�v�K��P����
]�U�츈 �OV�>� u� ǆx�  ��x��B� ��x���x�� r�ǆx�  �.��z�Ğz�&�? t��~�&8w�&8Gr⋶x��B�D��x���x��F9�x�s��x��v� ��~�������z���|�밋v���Dt�ދv�F8 u� �+�^��]�U��. �aN�F� H�F� �F�P�F�P�c���F։F��F�e�F����F� �F����F�  �F�F��F�P�F�P�F�P�c��+�P�F�P�b���F�+��F��F��F��F�F��F��F��^�F��^�&�&�W������+�P�F�P��a����]ÐU�츪�MǆV�A ǆ�� ǆ�� ǆZ� ǆ�� ǆ��$ �F�� �Ɔ�:Ɔ� �v�� �P�?a���� �P�c���u�v����P�ba���F*�-@ ����P�� P��V�P�;6��J��t �� P+�PP� P� P����
� P�����F�F��F�:�F� �� P�ca��= t��P�F�P�`���� P�F�P�`���F�P�� P��`���F��X�ƆY�:ƆZ� � P� P�� P�����u�����P��X�P�[`����X�P��b���t �� P+�PP� P� P�����
�P�a����F����Ɔ��:Ɔ�� ��P����P�`��ƆD� ����P����P��Z�� P��������P+�PP� 6�ǆ�� ����� P��������P�36��J��t �� P+�PP� P� P�J���
�P������ % ��J�= t���P� P��_���u+�P� P�� P����V�>! .uW�>" 0|P�>" 9I�># 0|B�># 9;�>$ 0|4�>$ 9-�>%  u&� P� P�� P��������P+�PP�����ƆD���D� uMǆ�� ����� P��������P�36��J��t �� P+�PP� P� P�n���
�P������ u���D� u�"�������6��J�� �	��% ���T�� ���% ����� % �� �+ұ�ja����+����T�щ���������� �4�
�
�� P+�P� PP� P�����
����P�V���� PP�� P�����u����P�F*�P�F�P��L�P���� ����P����P�F*�P�F�P��0�P����� PP�� P�N����uE�v�v�v�v
�v����P���������F*�P�FP��\�P��0�P��L�P��~�P�F�P�f�E�v����P�v�v
�v������������P�F*�P�FP��\�P��0�P��L�P��~�P�F�P���"��P�L��� P�@ P�� P�����~��u�� P� P�� P�����t-� P� P�� P�p���= t� PP�� P�\����t�� �>��t�6��6��������+ҹ
 ��0��V�����+����0��W�ƆX� �F��F�ƆG� ��V���� ���V�P�]������F��	����F�P��\������ P+�P� PP� P�����
�� P� P+�P� P�
 P����
ǆ"�D�� ,@��$���"�P��"�P�V]�������]�U��x �HV�F� �F����F� �F� �F�$ �F
�F��F�:�F� ��P�F�P�[���F����F� �F�P�F�P�v�� P�v��F�P+�PP� 6�F��tc�� P+�PP� P� P�	���
�P�����O�F� �v޸ P�v��F�P�36�F��t �� P+�PP� P� P�����
�P�H���� % �F�= t��vޚ�6�F��>" .u1�># 0|*�># 9#�>$ 0|�>$ 9�>% 0|�>% 9�>&  t �� P+�PP� P� P�U���
�P������~� t� �^�F�9t+�P�@ P�� P����F� �F
�F��F�:�F� � P�F�P�]Z���F�P��P�F�P+�PPP� P�� P+�PP�!6�F��t �� P+�PP� P� P�����
�P�F����F�P�� P��P�6��\��
�F��uo�F�+�=� ue� �
�.$ �Ȱd�.# ��Ƞ% �ȁ���N܋^��9u�B��� P+�PP� P� P�N���
�� P� P+�P� P�
 P�5���
�F�  ���� P+�PP� P� P����
�P������F�^�^�v&�D	�G�^�v&��� ��F
�F��F� �F���� ��F�P�Y����� P� P�� P����u�� P+�P� PP�  ��� P+�P� PP� P����
� P� P�� P�W��= uW�^�G*�
��0�F�G*����0�f��F� �F��� ��F�P�'Y������ P+�P� PP� P����
�^�v�D*�@�^��]�U��" �~DV�F� �F�F��F�:�F� ��P�F�P�/X���F�P�F�P�F�P+�PPP� P�� P+�PP�!6�F��t �� P+�PP� P� P���
�P����F�P� P�v�v��vZ��
�F��u�~�} �� P+�PP� P� P�T��
�P�����^�
�gG�^�G�^�g*��O*���F��^�v���v��6�~� uu�^�G*�^
;t+�P�@ P�� P�����F� �F�F��F� �F���� ��F�P�W����� P� P�� P����uW�� P+�P� PP�  �U�^�G*�^
;t��� P+�PP� P� P�u��
�� P� P+�P� P�
 P�\��
�F�  �`��� P+�P� PP� P�>��
� P� P�� P���= uW�^�G*�
��0�F�G*����0�f��F� �F���� ��F�P��V������ P+�P� PP� P����
�^
�v�D*�@�^��]ÐU���7BV�F� ǆ<�  �F�  �F����F� �F�$ �F��H�ƆI�:ƆJ� �v��H�P��U����P��H�P�U����H�P�F�P� P� P�v��F�P+�PP� 6�F��t�n� % �F�= u����P� P��U���u���~�u�6��6��F� � P��>�P�U���v�v�v"�F*�P�FP�v��6 �6 �6 �6 �6 ��>�P�v����F��t�o� P� P�� P�|��= ux��P�v�NU���u�D��P�v�:U���u�0��P�v�&U���u��P�v�U���u��P�v��T���u���P�v��T���u��� P�  P�� P����= t9� P�  P�� P�����t��v$�F*�P�FP�v�K���F��t�� P�@ P�� P����u��<� u�^�Qt�g�^�Qu�F�9GQt �� P+�PP� P� P�z���
�P�����F P����P��S���F P�FT��= t�P����P�S���v����P�S������P�T���F���Ƃ���v�Ƃ��
�v�Ƃ�� �F� @�F� ����P��S���F����F��F�P�F�P�T��� P� P�� P����u+�P� P�� P����?�F�P�v�v"�v�v�F*�P�FP�v�v
�v�v�v�F�P�v�v�v�v���"ǆ<� � P� P�� P�B���u� P� P�� P�,���~��t-�F�  ��F� �v�� P�v��F�P�36�F��~� u����6��6�~�t�~� t�v��@���v��f���~��t�v���6�F��tP����v��A��^��]ÐU�� �=>�F�F��F�F��

�tF�F��F��^���F��^�8t� PP�� P�h���u"�^��? u�^��?\t�^�?\u
� u+��� ��]�U�� ��=�F�F��F�F��^��?*uo��F��^���F�<.t
�u�? u$��F��^���F�<.t
�u�? t�.u0+��k�^��*u���F��^���F�<.t
�u�? u)�^�� tи �:�^���F��^�8t<?u�^��? t��F��F��e��^��?.uπ*uɋ^��? 돋�]�U�츈 �=ǆ|� ǆx����F� �F� �F�$ � P� P�� P�;���uq�^�GW�	��% ��F��GW���% �FҋGW% �F�P�v��v�� P��?���^
�w"�w �w�QP��?���^
�F�9Gu�F�9G u�F�9G"t� �� PP�� P����u9�^�GU���% �F��GU���%? �F΋GU% �F�^
�F�9Gu��F�9Gu��F��~�Ɔ�:�F� �F P��~�P��O���F P�[P��= t��P��~�P�O���v��~�P�O����~�P�F�P��z�P+�PPP� P�� P+�PP�!6�F��t+�P� P�� P����+����v�� P�F�P��|��	6�F��tP�'���v��M����~�P�F�P+�PP�Y6�F��tP�����v��"���v��6� P�� P�� P�t���u��� P� P�� P�[���t� P� P�� P�E���u&�F�	��% ��F��F���% �FҋF�% �Fظ P� P�� P�	���u6�^
�F�9Gs�+�u�F�9Gs���F�9Gu�F�9Gu�F�9Gs��� P� P�� P����u6�^
�F�9Gv���u�F�9Gv����F�9Gu�F�9Gu�F�9Gv��� P� P�� P�q���t� P�  P�� P�[���u#�F���% �F��F���%? �F΋F�% �F� P� P�� P�"���u4�^
�F�9s�E�u�F�9Gs�8��F�9u�F�9Gu�F�9Gs��� P�  P�� P�����u6�^
�F�9Gv���u�F�9Gv����F�9Gu�F�9Gu�F�9Gv���� P�@ P�� P����u�F�%  �F�=  t��� P� P�� P�e���t�t��F�% �F�= t�F�%  �F�=  t�U��F P�v�F*�P�v������F�= u�O��.���]�U��� �8�^��F��v�hP�L���F�F��F�:�F� �v�F�P�ML���F�P��P��6�P+�PPP� P�� P+�PP�!6�F��t�� P+�PP� P� P���
�v��#����z�P�� P�P�6��N��
�F��t�� P+�PP� P� P�u��
�v�������z�� t� �� �
�&�*���^�GQ�>!\t�>!/uظ!P�F�P��K����|�P�F�P�F�P��8�P�F�P�M��
��8�P�v�E���= t��|�P�v����= u�^�F���}��^�F
�GU�^�F�GW�^�F�GS�^�F�V�GY�W[��|�P�v�@K����8�P�F P�.K���>�u	�^�GP��^�GP �^�F��+���]�U��t ��6+��F��F��F��� �P�@K�����F% �F�= u�� P�� P� P� P� ��� P�� P� P� P� P���
�F�#e�u�F��F�P�F�P�! P�*K���� P+�PP� P� P����
�~�w��~�ur�F�F��F�:�F� �v
�F�P�J���v
�J��= t��P�F�P��I���v�F�P��I���F�P+�P�v��v���6�F��tP����v�����+��� ��]�U��� ��5V�F� �F�  �F� �F�  ��	 �F�P��P�F�P�F�P�v �v��	P�F�P�v�k���F��t�=�^�H�FފF�F��F�:�F� ��P�F�P�-I���F�+ҹd ��0�F�F�+���Vދ�+ҹ
 ��0�F�F�+���VފF�0�F��F� �F�P��P�F�P+�PPP� P�� P+�PP�!6�F��t�� P+�PP� P� P�W��
�v�������P�v�
I���tU��P�v��H���tD��P�v��H���t3��P�v��H���t"��P�v��H���t��P�v�H���u��P�F P�H���u��� P�  P�� P����= t9� P�  P�� P�����t��v$�F*�P�FP�v�����F��t�|� P�@ P�� P�S����u�~� u�^�F�9GQt�R�^�F�9GQt �� P+�PP� P� P�5��
�P����F P��:�P�G���F P�H��= t��P��:�P�OG���v��:�P�AG����:�P��G���Fԋ�Ƃ:��v�Ƃ;�
�v�Ƃ<� �F� @�F� ��:�P�G���F�:��F��F�P�F�P�UH��� P� P�� P�k߃��u+�P� P�� P�V߃��>�F�P�v�v �v�v�F*�P�FP�v�v
�v�v�v�v"�v�v�v�v����"�F� � P� P�� P��ރ��u� P� P�� P��ރ��>�	u6�F� �F�P��P�F�P�F�P�v �v��	P�F�P�v����F��u�y��6��6^��]ÐU��X �32V��F��^��0"�����^�?ud�^�?u\�F�\�F�  �v��^�&�@�B��F��~�?v��F� �F�P�v
���= u�^�&�B�uM&�D�uF�^� �^�  �^�? uU�^�? t����P�v��E���t�� �F�P�F P�E�� ���F�\�F�  �v��^�&�@�B��F��~�?v��n��^�T��>�u���&�G*�% �F�= t:�^�? t��^�? u��^�&�B�u&�D�u�^� �^�  ����[����F�  �v���&�@�B��F��~�v��F� �F�P�v�����u��^뽋^�G\�^�G �v�F P�|D���F�  �v���&�@�ދv� �F��~�v�^�G �^�6�&�D�GP�^�6�&�D�GQ�^�6�&�D�GU�^�6�&�D �GW�^�6�&�D�GS�^�6�&�D&�T�GY�W[�^�6�&�D&�T�G]�W_�^�? t��^�? u.�^�&�B�u&�D�u	�^�  ��>��^�v�&�D@����^�F��V���W�^������W+��� ^��]�U��Z �/V�^��W�F��V��^��W������P�v�C���F�\�F�  �v��^�&�@�B��F��~�?v��F� �F�P�v
������t�� ��&�G*�% �F�= t=�^�? t��^�? t� �^�&�B�u&�D�u�^� �^�  � �G� �F�  �v���&�@�B��F��~�v��F� �F�P�v������u/�^�  �F�  �v��^�&�@�ދv� �F��~�?v�^�G? �"�^�? t��^�? u�c��6�3��^� �^�F��V���W�^������W�v�v�v�v�v�v
�v�v�v������F�^��]�U�� �.��P�v�B����F��^��� �>�u��^� �^� �^�F��V���W�^������W�v�v�v�v�v�v
�v�v�v�p��F���]�U�� �-�6��6X�6V+�P�F�P��6�F��F�P�F P�P�6���C��
�F��t �� P+�PP� P� P��݃�
�P�7܃����W ��]�U�� �--�F�P�F P�P�6��C��
�F��t �� P+�PP� P� P�u݃�
�P��ۃ���� ��]�U�� ��,�6�+�PP� P�F�P��6�F��t �� P+�PP� P� P�#݃�
�P�ۃ��F�P� P�ZP�6��C��
�F��u�~�t �� P+�PP� P� P��܃�
�P�Nۃ��6��v��v�+�P�F�P��6�F���]�U�� �2,�F�P�Z*�P�0"P�6��B��
�F��t �� P+�PP� P� P�x܃�
�P��ڃ��� �0"������]ÐU��N��+V�F�  �F� ǆr� ǆn�$ �F� ǆh� �F��	��	:��	 �v��	P�i?���F*�P�v����F�= u�� P+�PP� P� P��ۃ�
�u+�P�� P�� P�׃��^�GY�W[�F��V�� PP�� P�׃��u	�n�� �^� �v
�v�v��v���A�������v
�v�v��v��BB��~��V��u�t
������ ǆv� ǆx�  �� �v
�v��v���x�- �� RP�_A�^G]W_��j���l��6�RP+�P�F�P��6�F�������9�v�u'9�x�u!�v
�v- �� RP�A)F�V���f�P�v����f�P�v�6^�6\�6���@��
�F��6��6^�6\��f���p�P��6�F���p�9�f�t�F*�P�v
�v�m
����v���x� ������9�x�wUr9�v�wM� PP�� P�Bփ��t�����f�P�v�6^�6\�6��;@��
�F��u�l�P�uڃ��v��؃��Y��P�v��=���tU�P�v��=���tD�P�v�=���t3�*P�v�=���t"�1P�v�=���t�;P�v�=���u+�P� P�� P�Ճ�� P� P�FP P�xՃ��t� �F*�P�v���� P� P�� P�PՃ��t��� PP�� P�:Ճ��t���F���Ɔ�:Ɔ� �v���P�<���OP���P�w<���F������P�F�P� P� P��n���r�P+�PP� 6�F��u���\� PP�� P�ԃ��u'�6��6�~� u0�^$��F��F� P��6�F���6��6�6��6�����>��t�6��6�����CP�L+���^"�+ҹ
 ��0�F��+����0�V��F� �F�F��F� �F���� ��F�P�&<�����F��	���F�P�<������ P+�P� PP� P��׃�
�� P� P+�P� P�
 P��׃�
�F�D�F�F�F�P�F�P�<��� PP�� P�Ӄ��u�v"�F*�P�v�v�����v�v"�F*�P�v�v�v��ރ��F�� PP�� P�RӃ��t�E�F���Ɔ�:Ɔ� �hP���P�:��ǆt������P��t�P�v�� P��n���r�P+�PP� 6�ǆr� ��t�� P��n���r�P�36�F��t�� P+�PP� P� P��փ�
�v��LՃ�� % �F�= t���t���6�F�� P���P�A:���v"�v�v �F*�P�FP�v��6 �6 �6 �6 �6 ���P�v�F���F��t�� P+�PP� P� P�Uփ�
�v���ԃ��^�F�9GQu�N�� P+�PP� P� P�(փ�
�P�+�F�P��P��z�P�F�P�v�F P��	P��h�P�v�Z����F�� �� P+�PP� P� P��Ճ�
�P�Hԃ��~� uڋ^�F�9GQt �� P+�PP� P� P�Ճ�
�P�ԃ��^"�H�F��F�F��F�:�F� �EP�F�P��8���F�+ҹd ��0�F�F�+���V���+ҹ
 ��0�F�F�+���V��F�0�F��F� �F�P��P���P+�PPP� P�� P+�PP�!6�F��t�� P+�PP� P� P��ԃ�
�v��iӃ�+�P� P�� P��Ѓ��F P����P�d8���F P�8��= t�MP����P�8���v����P��7������P�8����|���Ƃ����|�Ƃ��
��|�Ƃ�� �F� @�F� ����P�V8���F썆���F�F�P�F�P�9���u�ǆr� �v�� P��n���r�P�36�F��t�F���� % �F�= tɸRP� P��7���t�hP� P�7���ue�v�� P��n���r�P�36�F��uB�_P� P�7���t�hP� P�v7���u#�v�� P��n���r�P�36�F��t�F����^$�F��+�P� P�� P�Rσ�^��]�U�츞 ��"�F����F� �F� �F�$ �Fa P�F P� 7���tj�F P�Fa P�6���F��b�Ɔc�:Ɔd� �Fa P��b�P�S6����b�P�8���t$�^�GP*�P�FP�� P�S ���>� t+��A�^�GP*�P�h���F��t��	P+�PPP��6�F��^�GP*�P�@���F��t�� ��]�U��t ��!V�F� �F�F��F�:�F� �v�F�P�5���F�P�F6���F��F����`�~� uh��N��v��z�\t7�}�� P+�PP� P� P�҃�
�� P� P+�P� P�
 P� ҃�
�F��v��B� �F��v���F��B��F�P�7���u��F��F��~� |S�~� uM�v���r��B�\�F�P�t7���tN�� P+�PP� P� P�у�
�� P� P+�P� P�
 P�~у�
�F��F�P�:7���F*�P� ���F���N��^��]�U�� �� �F�  �F� l�F� �F� �F�  �F��F��	�F����F�P�F�P��5���F�t�F��F��F��F���]�U�� �x �F� �F*�-@ �F��6�� P�F�P� P�	6�F��t�� P+�PP� P� P�Ѓ�
�v��4σ��^�GW�F�GU�F��6�� P�F�P�v��6�F��t�� P+�PP� P� P�gЃ�
�v���΃��6��6�^�gS߸�	P�^�wS+�PP��6�F�� P�� P�� P�
�+���]�U��
 ��F*�-@ �F�P� P�v�� P��6�F��^��w�w�w�w+�P�w�6RP��5�F��V��F�V9V�wyr9F�sr�� P+�PP� P� P�σ�
�6��6��	P+�PP��6�F��t#��	P+�PPP��6�F���	P+�PP��6�F��� P+�PP� P� P�Wσ�
�p ��� P+�PP� P� P�<σ�
�P��+���]Ð�y  ��&�6��l�n  ��  �r  �>[]�@|<�B>+�D=;�gs���S&�&:s� [��6{SWU���z u>���r7�[t2�u�z u�&�"�zAtN��<=u�zC��sɬ�C��N�6p� �&��6��</t1�<"t�zuP&�G2�9ls�l��CC�&�� �f�n �^&�G2�@���&�2��tCS&�� [s?CC���n �3&�G2�@���&�2���@�&�2��tCS&��T [s
CC���n ]_[�l�n�6p�r�t��P&�� u�l�< u� u�n �P���� X��X���UQ&�O2��t�o	�\s� �����.��Y]�&�~  tE��EÀz���rB�&z�P�}+�{X�6}�< u#�|�:u�n	 �&�? t&� u�n �	� ����
P���� X��W&��>r&�&�eP��&�EX<u
&�U&�M�Y<u&�U�O<t�<t�<u&�U�=<u�{@&�E&�]�+&�u&�]P&�Gt��	&�Gt��� X&�Gt� _��G P&��uPSRW�n	 ����`�_Z[X�,� t�n  ���>n	u� t�n  ���>n	u��<�� t�n  ���c�>n	u#� t�n  ���>n	u�  t	�n  � �>Gu�>n u�n	 X�PV�
�t<:u�| u� �	�+sFF��^X�VR�Њ�r
�t� ��FF��Z^�<�s<arB<zw>$��:SW�>9��t�>48tPQR�e�»��� ����!ZYX�]�ECC,�&�_[�<0r<9w,0����PSRW&�&�
�u����n	 ����!�_Z[X�PURV���|r:�r��zt<=u&�~ un��zt<:u
&�~  uZF�Z&:F u
�tPFE�&:F uCF�E&:F u9FE��z@t&�G  t&�~  t"&� t<:u	&�~  u�< u&�~ :t���6}�^Z]X�PQRVSV� ^�,  �.  �0  � r�,
�t� re�.
�t� rY�0
�uR�
��t�,
�uB�ȡ.
�u9��0��u����,�.
�u�ȡ0
�u���ds��l[^�������[^�������n	 ZYXÍ6
�<�t�RP� 8���!XZ�QR3Ɋ
�t;�>	 t��u<:t0<.t,�<-t&</t"<.t�A�r� ��
 ���u�r�F뿊���F�����ZY�PQRVSV���D^u�� �,  �.  �0  �2  �	��w�rS�,
�tU�k�rG�.
�tI��]�r9�0
�u/�yu4�6p�|�,u*�D�.�y  �y��&�6����"�rX�2
�uQ�,
�uJ�yt<w?u2��zt<tr,<w(�С.
�u��0
�u�ȡ2
�u��[^������[^����~��n	 �	 ZYX�PV�F
�u��D� <pt<at<mu N�D� <pt<at	��z��y�D� ^X�PWV�>{�
�t�W u �G^� _�9^� _&� u-�n �%XV�
�t�* t�[sGFGF��t� G�>p^_X� t	P������X�SQ�>�	 :tC��AY[�PR�
�t5�r*�|:t&� t�| u <ar<zw,`�д������n	 ZXì�  t�Q u�z t��zAt	N����N���SQ<t-< t)<
t%&�}r3�&�]��&�9 t3�&�	C&:t��<Y[�SQ�t �&z�< t6<	t2<,t1< u�< u� F:��&�}r3�&�M�t� C&:t��< Y[ât�zu�z :���.�;�t</u�P�G��^�r��W�X���
</u�z@��VS�>w u%PQRWU3��޸ c�!���]_ZYXt%�6u�w�6u�w�< t:r:Dw��FF���[^�U��WV�~�E
P��]�M�U�u_U��]W�~��]�M�U�u��ĉEX�E
^_��]�PSRW3Ɏ�3��.� �/6�R6�>P�.��/6�Z6�>X�.��/6�j6�>h�.��/6�N6�>L��e  6�J6�>H6�f6�>d�f  6�^6�>\�.��/6�r6�>p6��
6��$6��  6��
 ��e  6�v6�>t� �0 �C Q�R rY_Z[X�����PV� c�!r
6�6|6�~^Xø D�  3��!�����D�!ø D� 3��!���D�!ô0�!=u��= s����� � �  � ����PSQUWR��6��6�6��Y  �t#�u�/ ���rZ�_
�t�������_Z�r]Y[�������PSR6�����u�, ��w s�Y�  �!2�������t;�t� ���rZ[X���u�&��!��� s&�U�!����t	&��!GIu���WPS���ٰ��u+�K��[X_�3��tO�@�׃�u(�!P&��Z Xs��@B�!�&�=u��������UQ����Y�!s�;�t;��u��]ø' � �À��t�ƀu�>�� ����W6�>|�t&�= �t&:r&:Ew�GG��_�6��3ۓ�6�6��6�6���	v��7���0RA�u�t<��u�|
,u6�6�A�$��u�|
,u6�6�A���u�|
,u6�6�A�3��3�3�6�6��3��t!�%� &8%u
&8et:�u&��K�sGGBIu�V���t5M6�>� u,�D0&:Eu�<0u�t4��6�>��uBBIIOO����W+����_Ys� Q�ʀ| t�tIIGG�^��u^�	���u3��tcUWQ3�6�>� u8�Du�|��%�Dt�Dt�Du�|���Du�g� ���" rY_]^���
�6�>� ur��6��  �3�6��6��
 �|�X6���C��@u���u�
6���CC���VS3�3ɀ��u	6ļt���(��t	6ļX���= r=' w	6ļd���6ļH�Ã��u���u��6������ 3����� t�T ���r�u뚜��u)RUQWP� �/<�Xu	�ظ�/��s_Y���� ]Z�����[^�WP���2����IX_Ã�u!6�>p�t=��uP6��6�pX�6�p�3ɀ��t&�M�	&85u&�M���s+��t���t&;�&;u�	It�����r
����u &}r2�&�G6�� �3ۀ| u6Ǉ� -CC6Ƈ� C� ]3�3�6���D	:�v*����D�t�D
6���C��@u� ��u�| t8Ls*L�ъL�t%�Du�Dt&�G�X6���C��@u�C ��u��D�u
�t�D
6���C��@u�$ ��u��Du�Dt�
�t	6����u�� U�QW��3ۍ>��.�r_Y�����]�D0u&�PA��s&�EP��&�
�tGA��+�U�]3�3�6�� 3��D u&&��Du��tC$6��
 �Du6��
 �X�Du(&��Du�ĀtC��6��
 �Du6��
 �*&�&�U�Du�ƀtC��6��
 �Du6��
 �D@t*PR�82����!s6��,�D
��ZX�D
,�g��ǈD
���\��t3Ҳ-RU�]6��
 �| 3�3�6�>� u � � 6�6�A3��D� 6�6�A�D�| 6�>�u �_ �n 6�6�A3��D�` 6�6�A�D�T 6�>�u�D�F 6�6�A�D�: 6�6�A� �. Uô8� ���!s6��  6��-ËD�Du=c v�c �6��6����I6:�u�0 PAA6�6��QR���v��$�������!��
�t�6�s�Ȋ��!����� rZY������+ �  �  �    * R	 y
 � �  " B g { � � �   ! H � � � � � �  �,	-I.�/�0�1;2v3�4�5H6�7�849p:�Incorrect DOS version
)
Source and target drives are the same
 
Invalid number of parameters
Invalid path

Invalid drive specification
+
WARNING! No files were found to restore
*
Insert backup diskette %1 in drive %2:
&
Insert restore target in drive %1:
!Press any key to continue . . .
L
WARNING! Diskette is out of sequence
Replace diskette or continue if OK
"
The last file was not restored
#
*** Files were backed up %1 ***
(
Source does not contain backup files

Insufficient memory
@
WARNING! File %1
is a read-only file
Replace the file (Y/N)?
Restore file sequence error

File creation error

Insufficient disk space
$
*** Not able to restore file ***
*
*** Restoring files from drive %1: ***
Q
WARNING! File %1
was changed after it was backed up
Replace the file (Y/N)?
Diskette: %1
Invalid date
Invalid time
No source drive specified
No target drive specified

&
*** Listing files on drive %1: ***
CRestores files that were backed up by using the BACKUP command.

QRESTORE drive1: drive2:[path[filename]] [/S] [/P] [/B:date] [/A:date] [/E:time]
  [/L:time] [/M] [/N] [/D]

F  drive1:  Specifies the drive on which the backup files are stored.
I  drive2:[path[filename]]
           Specifies the file(s) to restore.
>  /S       Restores files in all subdirectories in the path.
L  /P       Prompts before restoring read-only files or files changed since
A           the last backup (if appropriate attributes are set).
N  /B       Restores only files last changed on or before the specified date.
�  /A       Restores only files changed on or after the specified date.
  /E       Restores only files last changed at or earlier than the specified
           time.
M  /L       Restores only files changed at or later than the specified time.
?  /M       Restores only files changed since the last backup.
N  /N       Restores only files that no longer exist on the destination disk.
I  /D       Displays files on the backup disk that match specifications.
�>"]������ Extended Error %1�>�e�� ��� Parse Error %1�>f���U��WV�~�E
P��]�M�U�u_U��T  ]W�~��]�M�U�u��ĉEX�E
^_��]�U��WV�~�E
P��]�M�U�u_U��U  ]W�~��]�M�U�u��ĉEX�E
^_��]�U��3���F��]�U��3��V� �^*��6�� *�^��]�U��
 �eV+��F��F��>~u+�� � P����
� P������ P�F�P��P��	6�F��t�F��y�F�  �^��6
�F�� �^��6��F�� �F��~� |޸ P�F�P��P��	6�F��u����F��F�  �^��*��9v�t	�
�F�� �F��F��~� |��~ �I�^��]�U�� �V�F�  �v��怼� u��� u+��%�v���F8��w8��r� ��F��~�rǸ��^��]� �0�!<s� ���6 +��� r� ��ׁĞ"�s��3�P�v��L�!���6�&�6�&��Ʊ��H6����6 ��+��۴J�!6�������"+�3���; ��3��6�6�6肗P�� ���ظ 6��tiP�{���� P���0�!��� 5�!����� %��h�!���.��&�6, ����3�6��s�M6���ڻ 6����&�, �6��3�&�= t,� ���t��3��u����� ������tH���� �� �� D�!r
�t�� @Ky羦��� ����� �U�쾨���} �����t �U�쾨���f �����l � �t�~ u�F� � � �� t�>�!C��� �F�L�!���� ����� %�!�>" t�#�$�%�!�;�s
OO��������;�s���Et����� U��� P�{�>( t�(�� P�i��]ø �[�Y��+�r
;*r����3��E�V3��B 2���2�����Ut��� P�,� ^Ï,� 8�t)��&�, �3��� �3��u�GG�>�����ыѿ �� ���< t�<	t�<to
�tkGN�< t�<	t�<t\
�tX<"t$<\tB��3�A�<\t�<"t��Ӌ���Ѩu��N�<t+
�t'<"t�<\tB��3�A�<\t�<"t��ۋ���Ѩu���>�G��׀��+�ģ���6�?CC�6��
�u��� 6���3���< t�<	t�<u� 
�u�y�6�?CCN�< t�<	t�<tb
�t^<"t'<\t���3�A�<\t�<"t�\��Ѱ\���s�"���N�<t.
�t*<"t�<\t���3�A�<\t�<"t�\��ٰ\���s��"���3���  �&,U��U��3ɋ����I�6, �t��&�>   t�E�u�E�@$������W�	 � _�ϋ���.��3�I��<;Ct�~ EE��
�u���N ]��]�U��VW�V���;�t@�t�3��������_^��]� U��W�v����t���3�������I� �@�!_��]� ���r59�s% P�ر��ً�+���ËشJ�!Xr$�H����.��Ë���r3���]�s�P� X��]�s� ������]�2�� â�
�u#�>�r<"s< r���<v��.ט��Ê���U���WV�D+����D�tV�0��@tG��96\s��^_��]�U���WV�L�F�F�V�������FP�vV�a���F�VW�R���F�^_��]�U���WV�v�D��F���-D������������F��D�t�D@t�L ������Du�L�d�+��D���~��Du_�ށ�D�������������uF��Lt��Tu3�v�����u-�B��Lu�

���0 �D��^��G ���V� ���Du�ށ�D�������������tP�<+|�D@��^��GH�D�~W�t�v�����F����^���  t� P+�PPS��
���\�F���� ��P�FP�v��P���F�9~�t����F*�^_��]ÐU���V�F-D������������F�� P�\���^�G�t�O�^��G ���^�O�F�@�G�^��G �^��D��G  ^��]�U���V�v�B��Lu�F�

����Tu$�F�0 �Du�ށ�D�������������t+��5��-D������������F��F��D��^�� �G�D��L� ^��]�U���V�~ t[�~Lt�~Tuv�^�G�P����td�F-D������������F��v�K ���^�� �G  �^��+���G�*��^�

t�0 u�G�P�A���t	�v� ��^��]�U���WV�v+��D$<uF�Du�ށ�D�������������t'�+D�F��~P�t�D�P�c	��;F�t�L ����D��D  ��^_��]�U��d�!�WV�v�������F���F����  ��  �|�<%t�X�� +���������������������  �|0u<F��0 �3�<+u����  �"��< u�>� u������	�<-u���F��P�����u�V��P�f�����>� }�����أ��<.u#��FV��P�<�����>� }
�� ����=F t2=N t5=h t =l u�� �>� u�<LuF�< u��� ���� ���� �ӊ�����=E t
=G t=X u	������ ����-c = v���.���s���������i�����  �
 P����Q�� �������>� u	�� ����  ���� �>�u� +����F�9�t'���F��>� t	��  ���.����}+������ P�� ���: P�����~� t"�>� t�F�- ���}+�������  �.�� P� ����� �/�+�P���*��� ����������>� t��N��G�= t�=%u���+�PV�������< t�|��>� uY���G tO����M�s�r�s�s�s�s�r�s�s�s�s�r�r�r�s�s�s�s�r�s�s�s�>� t�>� u���G u��F뙐��^_��]ÐU���WV�~
t���>�t�>�u����W�F��V����*�>� t����F��F�  �������F��V����>� t�F�F�t�F�+����6��>� u*�~� }$�~
u�-F�F��V��؃� �ډF��V��F� ��F�  �F���vW�v��v���	���>� t!W�	����+ȉN����0F��I���N�����t<a|�, FG�}� u�>� u���t�~� u� �+�P���^_��]ÐU���WV�~ t� ���F��^���� �>�u����W�F��V���������F��F��^����>�u�F�F�u�^�	�~� u	�e�F��^��F��V��F�V�+�96�t�����^��F�&�? tF;�~��F�^��F�&�? u�>�+��>� uW���V�v��v��o���>� tW���^_��]�U������F��~gt�~Gu��*��F��>� u�� �~� t�>� u�� �6��6��v�6��v�����
�~� t�>� u�6������>� t�>� u�6���������  ���t�v������t� �+�P���]�U��V�>� u/���Ox�F�7��*���S�v����@u������^]ÐU���WV�>� uI�v�~B��6��6��]���@u����N�~���Ox۠��?��*��܃>� u�F�^_��]�U���WV�v�>� uP��6��^&��P�����@u���F��N�t���Ox��^&����?��*��҃>� u�F�^_��]�U���
WV�6�+��F��F��>�0u9�t9�t9�u��  �>�V�a���F�+�+~�>� u�<-u�>�0u��P�����N��>�0t�~�>� t�~ t�F��_ �>� t�F��j �>� u&W�����~ t	�~� u�5 �>� t	�~� u�= �v�V������>� t��  W�a���^_��]Ã>� t�+ ��  P����Ð�0 P������>�u�>� t�X ���x P�����ÐU���WV�v�F� �<*u���?��F�H��<-u�F���F+��<0|5�<909>�u�<0u��0 �����������ȃ�0��F�<0|�<9~�F�����^�?��^_��]ÐU���V�l�N��F�< t
:u�� ��+�^��]ÐU����^;�r� 	�*�F �tH�~
 t3ɋѸB�!rK�F
 uFVy(� ��6�V��F��ѸB�!FVy�N��V�� B�!�؋V�N�F
�B�!r�� ����U����^;�r� 	�����  t�B3ɋ��!r��� �tn�V3��F��F��WV����f��N�T�
�uJ�� =� vH���ܺ =(s�� +�ԋ��N�<
t;�t����# �a�;�u� ��
�F���� ��^_�U�E3���PSQ��+���^�@�!rF��tY[X��Ã�s�	��� @t�^�?u���� ��F�+F��f�^_���N�u�����V�@�!s�	���u��� @t
�ڀ?u����� ��Y�*;�s+�����3���U��^�t�O���]�U��VW�r�? u)� �su3���$@$��r�t�� ���D����6x�N�؎��	 _^��]��� At�������s�w�����tBH;�s���t4� ���D����t��L�+�H����L��ƌڌ�;�t&����&��=��t%���t��H;�s����t�� ���D���G�t���&��t�،�;�t&�|�7뼋w3��j ;�t$@@��^ t�M�� t�NN뙌،�;�t&����G3���Q�E��t+�IAA��&;�v��u����r�r��#�+�� u����u�3�Y�RQ� tW������D����w��+�J�U�XYZ�SP3�RRP� P� �����Z[t�� U��VW�~ u8���V�FHu�S r'�H�6�Ht;�t�D�FV�: ^s0�����s�u������ڃ��۱��H�!r钉�T�6�3�_^��]ËN��9Lt�����u���?��r9�ӎ�;�u9�s&����������;�u	١�+؎��J�!r;�u�������U��׋ތ؎��~3�����u��~������+����F�� t�I�������]� U��׋ދv���؎�3������ы~�Ǩt�I�������]�U��׋ތ؎��v�~3�������+��t������]� U��׌؎��~3�������I���]� U��VW� �HU��^;�}�� |�� @t� �3���]� U��VW��
�F�͋F�F�<%t
<&t�F����F���F�D�F�D�V�F��F�~��]�M�U�u�}
U�^�]�W�~��]�M�U�u�E
r3����� ��u��
_^��]�U��VW�~��]�M�U�u�}
�!W�~��]�M�U�u�E
r3���{� ��u_^��]� U��VW�~��]�M�U�u�u
�~��]_�!W�׎ߋ~��E�~��]�M�U�u�E
r3���� ��u_^��]� �N
�F�V�~W��
�t��
u�y
�-��ۃ� �ڋ��3��t�����0<9v'����u�O���D��D;�r�X_^��]� U��9�U��;�V�!�z�U��:�V�!s�= u쒓�C< t
<?t<*u�����U��?�U��@�^�N
�V�!r�^��7� U��F�^
؋^u�F���]� ��ȋF�f
ȋF��ы�]� 2��������� U��SV�F
�u�N�F3���؋F����8�ȋ^�V�F���������u�����f
��F���r;Vwr;FvN3Җ^[��]�  U��S�F
�u�N�F3���F���3��E�ȋ^�V�F���������u�����f
��f�r;Vwr;Fv+FV
+FV���؃� [��]� h� : e � � � < U��SQRVWU��ؾg� �~&�=��t= t#��� �u� �&��I� �t����� ��� �%�� �~&�5�/�!�
 � � � ��!�~
&��  &�  =  u�� �V�N� N�!s�� ��؋F� �~�> � �. #s� � �6 �> �D&�&�E&�E�D&�E&�E&�E
�D&�E&�E�D&�E&�E&�E�t&�e �&�E 3��D&�E� �  �@< t&�AC��&�A ��&�E��> � �~
&��  t� O�!r	�> �X�+�P��؀>  t�  �
 ��!X]_^ZY[��]� U��SQRVWU�^�V�N
�@�!r�v�+�]_^ZY[��]� U��SQRVWU�V
�A�!r+�]_^ZY[��]� U��SQRVWU��؋v��u�g� �u� ���$�3�]_^ZY[��]� U��SQRVWU���F
 �t+�v�<ar<{s�,Ar<s2�@@���v��� � �� �V� C�!s= tC� �N��v� �F% = t
= t= t2� � �v�  �V�F
�=�!r}�v��d��F% = t� �e��v� �V�N�<�!rQ�v��V���ظB�!r>�v��V+ɴ@�!r.�v��>�!r#�V�F
�=�!r�v���۸��؋F��� +���]_^ZY[��]� U��SQRVWU���ؾ �V�G�!r3�ߎǿ �� � �򮺀 +��~&�;�s� ����&��~
� �+�]_^ZY[��]�
  U��SQRVWU��!.����v
@����؍>� W� P+�P�x6�>�  t�����   ��   ��� ��� ��  � ��� �!��!2�;� t���ѝ� �� �>� |ٿ  �>� ~ϴ.���!��.� �� �� �v��\3�]_^ZY[��]� U��SQRVWU�V� C�!r	�v
�+��� ]_^ZY[��]� U��SQRVWU�V�N
�C�!r3�� ]_^ZY[��]�
 U��SQRVWU�V���F
�^�B�!r
�v��T+�]_^ZY[��]� U��SQRVWU�^�v�T�L
�W�!r+�]_^ZY[��]�
 U��SQRVWU�^����y� >�!r+�]_^ZY[��]� U��SQRVWU�^�� t������� t����������� �H�!r�v�+�]_^ZY[��]� U��SQRVWU�V�6�!=��u�W �r�P��P�� �� �� X�� �F<t�W �O��F= }�o �A��~+�&�&�E��+�&�E�� &����� &�+�&�E�� &�E+�&�E�� &�E+�]_^ZY[��]�
 U��SQRVWU��؋v��u�g� �u� �� �4����6 �/�!�
 � � � ��!�~&��  &�  =  u� �F
� �~�> � � O�!s� �. #s� � �6 �> �D&�&�E&�E�D&�E&�E&�E
�D&�E&�E�D&�E&�E&�E�t&�e �&�E 3��D&�E� �  �@< t&�AC��&�A ��&�E��> � �~&��  t�Y�+�P��؀>  t�  �
 ��!X]_^ZY[��]� U��SQRVWU�F=  ue�F=  |]= ?����=  ����M= 
������>= ��������-= 
������= t= � ���&���,��� �+��v
�]_^ZY[��]� �6�6U��SQRVWU�F= t� �<��F= t= t� �)��#5�!�v��D�V.�.��ʎںx�#%�!+�]_^ZY[��]� WVURQSP���؎�.�X[YZ]^_�WVURQSP���؎�.�X[YZ]^_���U��SQRVWU���ظ$5�!.��.���ʎں��$%�!3�]_^ZY[��]�     �.��<u�#�U��SQRVWU�^� W�!rp�v��L�T�L�T�L
�  �  �^�B�!rLRP�  �  �^�B�!�v�D�T��t	% � �� �D�TZY�^� B�!r���؋^ۋ� �F+�]_^ZY[��]�
 U��SQRVWU�v
��v�N�<ar	<{s��D���]_^ZY[��]�
 U��SQRVWU� c�!r�~�N�&�FG��3�]_^ZY[��]�

� _� � % �MS Run-Time Library - Copyright (c) 1988, Microsoft Corp9 � � ��    /B /A /Z /E /L /Y /S /P /M /N /D /? LPT1 LPT2 PRN CON NUL AUX LPT1: LPT2: PRN: CON: NUL: AUX: \ \*.* \ \ \ \ *.* LPT1 LPT2 PRN CON NUL AUX LPT1: LPT2: PRN: CON: NUL: AUX:   \ * * *.*  \ \BACKUP \ BACKUP*.??? BACKUPID.@@@ 
  CONTROL.??? ��BACKUPID.@@@  .* BACKUPID.@@@ IBMBIO.COM IBMDOS.COM COMMAND.COM MSDOS.SYS IO.SYS CMD.EXE \  ***DEBUG*** Restore file date is %02d-%02d-%02d
 ***DEBUG*** Requested date is    %02d-%02d-%02d
 \ \ BACKUP. IBMBIO.COM IBMDOS.COM CMD.EXE COMMAND.COM MSDOS.SYS IO.SYS \ \  no path from fnext no path from fnext no path from fnext  IBMBIO.COM IBMDOS.COM COMMAND.COM IO.SYS MSDOS.SYS CMD.EXE 
 BACKUP. \ .* BACKUPID.@@@ BACKUPID.@@@�� � ��� � ( ��    �    []|<>+=;" �  ����� �  ����� �  �� �    ����       
     
  �$A �MS DOS Version 6 (C)Copyright 1981-1994 Microsoft Corp Licensed Material - Property of Microsoft All rights reserved @(#)rctomid.c	5.1 86/05/13  B@(#)cmupper.c	1.1 86/06/17  `      �i  �� � L ��;C_FILE_INFO �  � ��� �  ��C �  ��#   	��                       �      B � x �   � t ��(null) (null) +- # �  �     @j@j@j@j@j �  �dm<<NMSG>>  R6000
- stack overflow
  R6003
- integer divide by 0
 	 R6009
- not enough space for environment
 � 
 � run-time error   R6002
- floating point not loaded
  R6001
- null pointer assignment
 � �� ��������������g    P�w	RB��� �  ��� ��O����P�4 PˌÌ�H�؎�� � ���G����H��� ��������+�s��+�����ڋ������+�s��+�����¬��N���F��$�<�u���<�um�¨t��2� �3ҭ�����Î�������t&��� �t�� �܌�@����&H����Ë> �6
 � - �؎��  ��֋����.�/�@� � �ʎں�!��L�!Packed file is corruptb � � z q X ^	f�v�D4�x�^v4X8`!�##�"�"�&&�+�+�(�(�+/ /�.�.�1N48L5>�=�<B�A�A@�?�ED�C�C;B%BB.G�F�F�J�JkJ<J�IHPK?K)KKUUZU VBf�fu��ńQ�|����+������n�r���%�ڌgg!gh�	h�h��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        MZ�     � ��� {)J�     � �U� �� j	                                                                                                                                                                                                                                                                                                                                                                                                                                                                              ���� � ) SETVERXX K        .� .� �S.� �G��u�����G[�PCMN 
KERNEL.EXE 
DOSOAD.SYS EXTDISK.SYS REDIR50.EXE 
REDIR5.EXE REDIRALL.EXE REDIRNP4.EXE 	EDLIN.EXE 
BACKUP.EXE 
ASSIGN.COM EXE2BIN.EXE JOIN.EXE RECOVER.EXE GRAFTABL.COM LMSETUP.EXE STACKER.COM 
NCACHE.EXE NCACHE2.EXE IBMCACHE.SYS XTRADRV.SYS 2XON.COM WINWORD.EXE
	EXCEL.EXE
LL3.EXE
REDIR4.EXE REDIR40.EXE MSREDIR.EXE 
WIN200.BIN(	METRO.EXE                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               SQ�0�!Y[=t3��3V�ȎؾK 3���t@@�����@^SP�R�!X�&�] K &�_ �[�G�O���                 U��R �mV��P�v�v�G�����|	V�J �����t:���؋��6�F�P����������F�P�����F�P�N���6<�D����^��]�U�� ��V�~u�@P� ��+�� �~u
�VP� ������ut�~u� ���g�~t�~u�?P�6�������}���`����u�~u����u+�S���u"�~t�68�����= u
�6:����u��~t���u��hP�
 ���^��]�U�� �1WV+��W�Y��F�^����؋?�u�^_��]�U��8 �V���F��F؉F��r� ��9F�r� �v��L���u����� �^���P��@P�F�P�����^������BȉF��	�^�� �F��F�9F�r�^���F��F��
 P�v��^��F���P�b���^���=
 }�s��vP�v������
 P+�P�v��Q��P�^��F���P�$���F�P�h
���^��? t�6���9F�u
�6>�K
��+�^��]�U��
 ����F��F�F���F��؊� �F���+�F��F�P�F��PS�a���F�F��F��v�+�P�v�����?P�v�� ���F��}�=��u'�0�F��t���N�+�+�P+�P�v��U��+�������]�U�� �hV�?P�n�������� �F��tC��+F�;�|9�^���,��?P�F�@P����^���@F��^��F��M��^��N�+�����^��]�U��3���V�=�^��P��@P�v�9���u�^���؋v�8 u	�F+��/�^�� F��9Fs�^�? tS� ���u��������^]�U��3��V�^������}�@;�s� �+�^]�U�� �c���F���^��� F��^��? t��;�r��;�s���+���]�U�� �&V�F�P+�P��P����t����� �F�P� P�TP�v����
�t� �~�t� �\���+�PR� P�6R�6P��P�v��U��
�ur� P�6p��P�����uW�>�uP����PR�6�������u����3�6��6R�6P�6��v��� ��
�u+���������������v������^��]�U��2 �(
V�F�P� P��P����t� +�P��P�����t� �F�P� P��P����ur+�P�6R�6P�v��%��;Pu,;Ru&�F�P�6��6��v��j��
�u��9F�u+������v��v��v��w���v������F�P��P�M��������^��]�U�� �_	+�P�v
�v�v���;Fu);V
u$�F�P�v�v�v����
�u�F9F�u+�������]�U�� �	WV�^�7�F@P�����~u� �8�F� ��^���~�1�I���F��F9F�|�xP�^�w�%���t�~~������ ���F� �: P�^�w����u� �^�_��-@ P����t|�^�_�:up�^�w�o���F�=C ~�����^�w�F@P����^��~�9\t�^�_� t�zP��@P����|P�F@P����F��F9F�|� �?����;�^���~�1����u��^��F���~�1�FE P����F9F�|����� ��P�^���~�1����t@�F��F9F�}/��P�^���~�1�����t�F��F9F�|X� � ���� � � ��P�^���~�1����t3�F��F9F�}7��P�^���~�1����t�F��F9F�}�����K�^���~��?/u����C�^��F���~�1�; ���F��t!�^�F��GS�^�F��GT�F9F�|�� ������������^_��]�U�� ��F�  �. P�v����F��tL��� �F��v�����F�= w�v�� ���u�F�����v�������
 �f��F��F��F�= r�0 P�v� ���F�~��tP�9��= w�v�8 ���u�F�  ��v�����*�	N��~�r�~� 
r�F�  �F���]�U��3�����^�F�������	u+���^�? u� ]�U��3����F�^�F8t��]�U�� ��^�F�?/u�^�? u+��&�^�F�8u�F�F�^��F�
�u�^�?��؋�]�U�� �J�. P�v����v�E���u� �v� ���u� �\ P�v����ut�v� ���ug�v�� ���uZ�. P�v�����F��t8�. P�F�@P�����u3�F�+F= (+�P�v����+F�H= � ��v�
��= v�+���]�U�� ��F� �^�? t�F��P� ���F��u�F���]�U�� �XWV�. P�v�L���F��t��� +�+����㋇��F��tP�v�M��= ��ً�G�tك~� t�^��.��^_��]�U��3����* P�v��
���u�? P�v��
���t� �+�]�U�� ���F�=  t=	 t= u�F�  �F��=/ t�=: |
=> ~�=| t��F� ����]�U�� �{+�P�v�r
���F���^��F8G�u�N��F9F�u�^�� ��]�U�� �A�F�F���F��P�f����u�^��?:u�F��^���F�
�u��N��F9F�r�^���F�<\t<:u��F��F���]�U��^���D�!s	= u3��� ]�U��V�v� ��
�t����!��	��^]�U���B�F
�^�V���!r�����]�VW�R�!S�0�!_��<~����ؾ	� ����tQWV��
�^_Yt	&�=��3��� _^� �0�!<s� ��6 +��� r� ��ׁ�n�s��3�P�v��L�!���6�&	6�&	�Ʊ��H6�	��6 ��+��۴J�!6��	����p+�3���; ��3��6�	�6�	�6�	�B�P�� ��ظ 6�	�P�{���� P�	�0�!��	� 5�!�s	�u	� %���!��
�.��	&�6, ��
��3�6��
s�M6��
�ڻ 6��
��	&�, �6��3�&�= t,� �f	�t��3��u������	������tH���� ���	�� D�!r
�t���	@Ky��
��
� ��
��
� �U������} ��
��
�t �U���
��
�f ��
��
�l � �t�~ u�F� � � ���	t�>�!C��� �F�L�!��
�� ��
�s	� %�!�>�	 t��	��	�%�!�;�s
OO��������;�s���Et����� U��� P�{�>�	 t��	�� P�i��]ø �[�Y��+�r
;�	r����3��E�V3��B 2���2�����Ut��� P�,� ^Ï�	� 8�	t)��	&�, ��	3��� �3��u�GG�>�	�����ыѿ �� ��	�< t�<	t�<to
�tkGN�< t�<	t�<t\
�tX<"t$<\tB��3�A�<\t�<"t��Ӌ���Ѩu��N�<t+
�t'<"t�<\tB��3�A�<\t�<"t��ۋ���Ѩu���>�	�G��׀��+�ģ�	���6�?CC�6�	��
�u��� 6��	�3���< t�<	t�<u� 
�u�y�6�?CCN�< t�<	t�<tb
�t^<"t'<\t���3�A�<\t�<"t�\��Ѱ\���s�"���N�<t.
�t*<"t�<\t���3�A�<\t�<"t�\��ٰ\���s��"���3���  �&�	U��U��	3ɋ����I�6, �t��&�>   t�E�u�E�@$������W�	 � _�ϋ���.�	��3�I��<;Ct�~ EE��
�u���N ]��]�U��VW�V��
�;�t@�t�3��������_^��]� U��W�v����t���3�������I� �@�!_��]� ��	r59	s% P�ر��ً�	+���ËشJ�!Xr$�H�	��.		Ë���r3���]�s�P� X��]�s� ������]�2�� â�	
�u#�>�	r<"s< r���<v���	ט�	Ê���U��^�t�O���]�U��VW��	�? u)� �su3���$@$���	��	�� ���D����6�	�N�؎��	 _^��]��� At�������s�w�����tBH;�s���t4� ���D����t��L�+�H����L��ƌڌ�;�t&��	��&��	=��t%���t��H;�s����t�� ���D���G�t���&��	t�،�;�t&��	�7뼋w3��j ;�t$@@��^ t�M�� t�NN뙌،�;�t&��	��G3���Q�E��t+�IAA��&;�	v��u����r�r��#�+�� u����u�3�Y�RQ� tW������D����w��+�J�U�XYZ�SP3�RRP� P� �����Z[t�� U��VW�~ u8�	�V�FHu�S r'�H�6d	Ht;�t�D�FV�: ^s0����d	s�u������ڃ��۱��H�!r钉�T�6d	3�_^��]ËN��9Lt����d	u���?��r9�ӎ�;�u9	s&����������;�u	١�	+؎��J�!r;�u�	�����U��׋ތ؎��~3�����u��~������+����F�� t�I�������]� U��׋ދv���؎�3������ы~�Ǩt�I�������]�U��׌؎��~3�������I���]� U��WV�~�v�ߋN��
�t���2���^_��]�U��WV�N�&�ً~��3����ˋ��v�D�3�:E�wtII�ы�^_��]��  U��WV�v3��3۬< t�<	t�P<-t<+u�<9w,0r���ҋˋ�����������؃� ��X<-�u�؃� ��^_]�U��VW��N�F3҃�
u��~� U��W�~��3�����A�يF���O8t3���_��]�U��֋v�^��
�t,��'C:�t�,A<ɀ� �A��,A<ɀ� �A:�t������]�U��^�ӊ
�t,a<sA�C�
�u�]�U��׋ތ؎��v�~�ǋN�*;�v���;�s����NO�����Ǩt�I�������]�U��׌؎��~�ߋN��F���� t�I�������]� �N
�F�V�~W��
�t��
u�y
�-��ۃ� �ڋ��3��t�����0<9v'����u�O���D��D;�r�X_^��]� U��^�>�!�a� U��O�V�U��N�V��!��Nu�V�N���!�8�U��V�F�=�!r�^��!� U��?�U��@�^�N
�V�!r�^���� U��V�N�C�!��� U��^�N�V�W�!���          MS Run-Time Library - Copyright (c) 1988, Microsoft Corp 
ERROR:  Invalid switch. Invalid filename. Insuffient memory. Invalid version number, format must be 2.11 - 9.99. Specified entry was not found in the version table. Could not find the file SETVER.EXE. Invalid drive specifier. Too many command line parameters. Missing parameter. Reading SETVER.EXE file. Version table is corrupt. The SETVER file in the specified path is not a compatible version. There is no more space in version table new entries. Writing SETVER.EXE file.An invalid path to SETVER.EXE was specified. 
Version table successfully updated The version change will take effect the next time you restart your system        Use "SETVER /?" for help 
No entries found in version table Sets the version number that MS-DOS reports to a program.
 Display current version table:  SETVER [drive:path] Add entry:                      SETVER [drive:path] filename n.nn Delete entry:                   SETVER [drive:path] filename /DELETE [/QUIET]
   [drive:path]    Specifies location of the SETVER.EXE file.   filename        Specifies the filename of the program.   n.nn            Specifies the MS-DOS version to be reported to the program.   /DELETE or /D   Deletes the version-table entry for the specified program.   /QUIET          Hides the message typically displayed during deletion of                   version-table entry. 
WARNING - Contact your software vendor for information about whether a specific program works with MS-DOS version 6.2. It is possible that Microsoft has not verified whether the program will successfully run if you use the SETVER command to change the program version number and version table. If you run the program after changing the version table in MS-DOS version 6.2, you may lose or corrupt data or introduce system instabilities. Microsoft is not responsible for any loss or damage, or for lost or corrupted data.  NOTE: SETVER device not loaded. To activate SETVER version reporting       you must load the SETVER.EXE device in your CONFIG.SYS. SETVERXX B L \ n � � � &H[t��Kp���:n� =v�\  ��W��*q  ���   .0 . ? \ SETVER.EXE DELETE QUIET QUIET DELETE AUX CLOCK$ COM1 COM2 COM3 COM4 CON LPT LPT1 LPT2 LPT3 LST NUL PRN  ��������������  
 SETVERXX     �                                                                              	;C_FILE_INFO                           ���                     �	C           p   	��                                (((((                  H����������������������                                                                                                                                                <<NMSG>>  R6000
- stack overflow
  R6003
- integer divide by 0
 	 R6009
- not enough space for environment
 � 
 � run-time error   R6002
- floating point not loaded
  R6001
- null pointer assignment
 ���                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 MZf�   V!��W    ��R   !PKLITE Copr. 1990-92 PKWARE Inc. All Rights Reserved   � �����|<`$� 0&                  ��?�O  ; r�	��!� Not enough memory$-  ��-% ���P�#3�W�D��ː���S��9 ڌ͋���������Ƌ���NN��+�+؎Ŏ�� ����u����� 3���� �8�����A����B����H����M����S����g����h����i���r���Jt�s�3�3���Jt�����Jt��Ӏ�s(��Jt��Ӆ�t��Jt��Ӏ�r��Jt��Ӏ�w}.��	��3ۃ�t*��Jt�r#��Jt�����Jt�����Ju����Ӏ�s.��/���V��+��^�u���Ju����Ӏ�r���Ju����Ӏ�r���Ju����Ӂ�� ��뻀���Ju����Ӏ�r��Ju����Ӏ�wE.����t�Z��Ȁ� <�s�M�P�� �����  ����Î��؋ރ���Î�X<�t)�������Ju����Ӏ�r��Ju�����.�����[���3�����Î���&����Ò���ҋ����S�P�Ŏ�3��؋ȋЋ�����      	
                    	
        U���
�F� �f��F  ��H�&�v�� `/�  k���r�4Q 0!<��آY �v
 � | ��
�u���=��>6� l@� P��0& �C��R �t%eJ�e�> u{	�c��&��6-�F���Ba:Wsaa��/u*��E��[ �q�;*  ���^&�w7L��!0���}t��I
 ^^�� �( +p#�ypOSڛ`x��H_6�H�G� �t� v���B P�v�u�2Q?��&�~�A9+��t�����R,E�+1N1l����t!�y6�J�z*l*��`J!f a�F��1��@�hu%�yd*��c�W�i�_��5u4��,�$��~(/(u����	��t*�����
�-�4@@9L� +�)(+�&����+H����v� ���]ːr|��Ȥ `N��M �n���&Ƈ���&Ǉ� ��]&���&������6��~��:P�+%���o��HR��.!9aT��3�VT�RX ��ZJH 8�l �j ��)��/���!JY����*�'� �] �g\��^�����{x����.�,�*��	x |��m�� ��������{O�V��tWV� T�!�~�� .^_���.�>�*3���333�X��r��
��G�X� [���?F=�D#+䠋�,� ����r,r�F+�*Pv�I �=�F��V�U�jz���~xL�:� �����J��F�AP]���9�=(�	��.~�	� �:�0	����>l� H���_Z9=��� u�<����T���Q�4A�h+�����~;;���R^�&��� ݉^���F�� 6�^�!G@Ո���?MWқZu TfR 9/w ��!
N�ON�7D� �����<��I����,��ߊԊ�*���,,f	�����F� �]M����Z�_��Rᇈ���9G��[��Un9	vr zf
}	�-R��  � Ɔgz�1�/�=��~�~��';��N�F�$ ���^P"^Q @&�� p��p���r��*�b��H=-t/��H ���� �	y�l���u$��'s�jw��!�,�*�Q�p=WE�)�)�(r)��N
8@A؉^��F �+u"��^Ȃ

0�HW2�x[3�.��`�x�����atĞI�y�SG�G[�#�� �t�� ��v����m�,&�,��^->>��נ� �m��808\'Qe�KT���vu3x����������S�5���]����v�u�����	��kf�
W7H�]�aݼ*�vuC�����%���>��U@ u� u5�,$	�� 9�������V��H�� e���uNT�@2�u�4�(��8��nK�� �� "r�4�����Վx/՗�զ?
lY�tZE�����VQ����U��*j����Z���d�� �����Hn3�>\�}l&�.I��d�Wr�}	��*wf��rY^dǆx�2�Y����Q���\
;��N�t��F����n���˛�Ly
��ŋ;A� 8��]H�
������uE��
�S�yZ�N(w��[�ѡ*]�]@�ɚ�&
�ٵ �4�@�D��M#� ,u#��&o��(T�P������<����+�P��+�QĠ�28�
`4�`5��d6�w6�7�Zv��(��7�F��+�^&8θGZv�����xo6�+'
�D��:0���&��-A �!c�Wq�<�d�z�&#hS�ɀ����:�0�t�b���A<�)� |��~�&�B���:�f�,���"�g��Ɂi�z�ucWI�Yt$���o�������#��`� /"�+/�,�kz�$
�� un�F8 Qt��&��P�#
��'u�
��V��ZDs|:��1�u6�"�,�\�<&L���a�e�����;uU��/R��L��� ��N�F&*<�t"�S+2+�Fȍ� ���jW���@�-77hZp�Vb+ �:Q�N
�VARQ�ܺ\ �2�FD�1�F@RP*�QR)'�Q�%I���*g@u(UJ�(�(���.+ Z��)+_�_���M���� �
���~�*��e8V�&f^~ �#9$=t��Y�}`؋v����� ��2��̐�� ,|H5rG���X�KG*�^� d�??��u��Ř�#\A
����0u\�}������l"T+t��Nst׾�բ�b��<ك�v
4,���qX� r)�(�(|�`�A%����p��t�@ꕒ ���
�EL
�
��
�
u��m�)R�e���H]�u��
]]

]�

-  �= w ���.���  $.8@HPXb�Tlv�Ǚ#��T�� �ڂ��� ������♙���֙����ʙ���������\R���&�  ��������@���0q� �ם/B#�V�Ip�$M#��P��]B���t$��$�3�^�����	��'$�W'I�(�&��u*t^a^��2f ��n~V�:�#��],������hh��yja N&��d�~�0D�zl%o�)V�<iv�r
["��~�C�T�6�M�K:!qn��>a"�W��Cw�]T��u�c��u�o�(z^�(&9M��ńΈ��w[\+�n�M7�{s�� �
��{�d��.���g�JpN=)^�r_I� ��+��骋��\Tt��`vb�Axg�Hlِ��C��.L��t諾����5�L_=�>��&
��&%hz�fx���|�:��N��к��3��{%�A๥���c�^7�64!��=�
k,~�ujc�$��b&����h�� ���t3�~�णz�:>W/Jk�f9"\� �]Q
p^V�|	FZ��*��i���i�0��-bCI�9u'Ǉ��v9j� j��"`�V/��EX.i�"�"6��)�"l�>�&n�g�}����̷�ÜuU�X�˅ S�ʶʶN�ʶ�ʶ��V#}���d����
���5��~�����@ ؀~�޵���h�$���,~��	�,q��{띐j.�\$9�����7��L��:�% @�������**/�5� �J��^-�� �~�h�Ў���J �?��S���X��s褀�� � -�y�� �8pA�P�x�NP)�Q���]FF��&V���MzKP{Z&%�&tD#�i_`&,�F�=�.���C���$��1^�{�������~��)��B��S�Fu��J�#���3dWw��g��`�&R@5�\�
�����Ɋʄ�u�T�;&;��@;�OJ*�����p4u8����/sP/~���$+�^�6�Z��#��S���O@.�3$Ⱥ�&^W녵����ۣ"��%�PRS��Bg��.ˢ�_RwN9	�S��~]L�骐�Ir��JR��[U{��%;� ��O��zҬg�y�Ɔ�� ���	 	P�NAQ��U@Q���i�~�jRZC(��|!r�� Q�O�
{�Rvw��i��4x����{��tyLn#tH��$�\TqЀ>�~X �u�'���4&l@p�6�������͚�2�\��P���Ū��~W%�#�rBI*u^K[�5!��ܣ-@���B�OOhz!@��o� ���E,��(�++�Z,��U��\��@\*�0a}���[=T�<�<�-hQ�yz(�|U��L*@�/���L��,�S�Ry�3D�WA6���6��5B����K�R�K2#?K7 �1���Z S��46&�haJ�,��F4Y6����i�_��]"f��� r������r"f�w>Q$�N�
@r�G8D�xF ���9��7�t.
�
����ֲ�`뉟�&D���DI�.
D����=�PI�@��T�qqc�U5��ty�Aq�qQ���⍿� ��;���B����C����5�'$(�aKb]\�y�d���U���2Jk����%��;P�����6��$�Lu!��6��X< [,ŽP	?��Wǆ��� ��� �Ƹ���u�ɼו�k�8]��q�2���0b�{	�	^�Fj�_E�iW��t�� �F
"�����5��g(P��P�l�P
��FP���8.CZD�A'���t "�H�����IR Huh)�@ua@@U	���T�_I��u
�PL�h���
c8�QW�':'-.fa)�,�j�,�e��b�l�F�D/��;W;"����	t�qTs�?��c� ��z�.V..g�%�%�٠ ۉ����d�5mu�J�Ru��c��`�@ؠ����ȱ"QU�
� a<�}?	aѭ�L�Ӷ=�g��f0�g��qhw:h��J h��h����h=4!Sw =�=z���E��
�U���
 ��nY?h0^!h�6�-!R^��ڱ�RUji'] i���i����F =��^=�� �	.)�|=]�Ԡ$
 c6]�c'�Vc�6R�N^^d'] ^���^��H�����j�_JQu!�YP��uw@J��@�!�Hu>t� �S���,�ҎFI���TY'�L������]d�i �C��*���^.e�����CF�e�0�e����@���~�U�tU�OS@�! �Sie e�7�f�EG:"!�� :�:�:�"��8b��<WVgp�F���F�=�g���њ�E�u=�5sd�V/~�L��aͥ����\�F��`��N���V̰NfJu �-  ���#�  �)�� ���#Ȁ��1futS�S�� ����^�W^��U�`����:�� �+j���#�K/	�N�q��L����y(��
� 3 �~� @w��"�������� ����뷢V�+��fH�	�7�	p���[1V&��� ��yf�)�)��`��#����x�NO��w>�*%Г�\���`���$��n���jg퐢t�9�d;� (�	a��{�u�P�M��7�$�t	�ȸ?�  ��!��Q�f��R�rT��&uQ�ݮ�F�t����ܚz,BHC�yp�dlf����������d.1�}�s}_�<Ou��--c�ut�$z7$�$L#RN $L*�:d��W#t'Qϓ�-H-J�I--7�0&3		��?��f���ц�,ίК�Qa$�N�pP�����������I���y�:);;7�N	7	 �c=��v+��s[;pr�]w;zv���Ћ`�_�f�ˋ���0&M�^/x�N� �+�;�w
r;�s�Ӌ��m��"��	uK����9F�u�	 L�@��ɐ��:0��	H���gt/�+�6�*4��*5��@���*5��5�5`���2��+�-�*�y9�U		ѓ�		� `<�u���'z���N�z�/!�'��+8I���{|o+0F�V���;V��r"��vI����`�V��T���}�� ]7=O���)�����2&�~�	�	u�wr�u�s�NFa�-���-���F��&!E�F!F�65
Eu/�����42[����`r�z��a��r�ڌ،ڴh���>�!�������/��f��I/�/�)����b��K}A{�}��0:F��V��=Y s�"`��v���e�en=ҋ����F���/��$j�lL�j%�L��>9�.p���-��(u�u��}u��m_�����&P�6f0!��e��:�&�k�u�R��6��T(�)U��5�u�BZ	/���ȐH=uv���~�9��*F�8T`W.	= Ts!	�Ԩd��iUس� �}5ࣘ�&���4 �1��&+*���pt:q7@��Y.��H<��5t �1�!�':c@�١l ���/��/�/�	 �0���)���/��/��A"u��on/M�/�/�$��D���ӟ�/�V鼚/�f�Nb��*�P/jJ�*/��,/~1$������/�Jꍖ�,/�	HQ�JB�J/[S/��/��x��N $��?-/L��I�/�$�" � �O�/5��/�1/'�H��Tb��/[S/��/�˸�)%$�褝�R��*JU�꥔w�"�h�fbhV�F� ڰ��^��������C. GU�,t�ݷ^�������,P*�I�~� |�y�E�%G&���G�� V�� WV�(�
���!�^$'U� AC��!�/�VdFV��
No w��t�+!Ʉ��|�����\
�N�kqBu<n)���u	 U���`��ݰ d��^ M�}������IF���f�����6�'-�-*�r�������)`V��Q��X�{�1���Ύ�Ht��/��D
��	�ڧ����D˸"}�/} �� C��MKNdK.T ���E��"4g `�'e' � �*2�&U��$��>��  J֔yp��
��L�Y��"��$ݼ�&m~N5��Dޘ*�(b�+�F��c J
���^��^��%Ü�r�q�^�>�~���1�$,]��TJ�%�r6��U]E�S����!��S��&�@��F�$<���W��.�ľ�f/�!.���uyVQ�v�tSN�B�TƇ� �z �_ J� Yt� x
 ��c0)�(Ҡ�* ��t   TPQRSTUVW�� �u2��!$ �_^][[ZYX� ϸ$��OK���x&p�(���ke6!�{�l��#�6(��)�!��i��x8�F�����J���/D��u= �V�.�Àt)��2��,�S��/�!x�[�^G������^��߫�c	����Qo�c��z/z ��`u`oS�
v�su;g@�9V�D�� !r�<�t2$����o������ ����zފHCI	��K��s�~Y��.�	.��D�/s+  Z+ +r�� ��t\1V��1�������3���
<	�7�$� �B: �^�9	�R,M�$�$ ��p��r,�;PU
3w j�9x���9�90�U9>�_9�9���99��^���~�0N���M�_�(�s>�N��	�_ �������S�X�V�|��hIUVW! |"��MDuB
 � O�7�N ��_^]�2��N�3���V�#Z#Z*��=�����(��<�T� te�Z Ƈ�������'3  ��A��g9L� h 2@���!^���<Il���*"�$	 [����,�#���d{�J^= ��Dܮ	L�D 3��F� ���^��^���~��3L�;�	�~]�s�]����@��F��]Ǉ��j��\��������z#�#��k#�#�}�#������kE=���f���N ��&�GH���ȴ�����+�+� �EH3,�8�P&��*%�=�����ө��� 0�WQ0�0שw��������p!����c`z�G*�W�6��R�l	�z�/Ͷ�/�f�S��<+�&�ѫ�����(��zg% ��= �'Jh���hP�� P��	H�w"
4@��Ƈ� m=f��ؽ6N�7�䋇@>�"�Ͱ�/w���7Ⱦ����G�� ls�;HF��V���h�Pԋ�� �DD�`�!s��z�8�ٖ�\�g���x����(��aqŖ�"@���</z�Go΢_��Ⅹ�!Ȓ������֫��\�x�鎆��'�0(K,0v���������R�m��K<Do�f�=N��H< -���7��H�7M��&?$��| ��&���E��f���@���hv�ʜ�~O�	�����7c��9�A���� Z\#w�Y�����Ym�^Q�R�H����������t�֍�F���1Bjhs�Dp����L����#�|��If��vN��`~�@s*L,��	�w>�� �+
Y� ^,W���X��E��  ES^� �w��s�y��@�Jer=�@� ��ꚤÄ�Y0� %���z���ǋ�*�)A������>�����������l�9Ft�$vM� ����ٸ g]� ��9Q�")��O ]��v;l*���~��X�#R�F}1�D�м{E�]�ƛ�$���@� ��zBK��LB;�H�U �z���}��P�dJP�JP@���
Ɔ~��W:��	H����-N���@P�3��4�N�TKg��ERz��� P|P
,���� ��g���`��Z`�G�W`��?	'1�!����r�+nj1rHQ��`b�Px QqN =}��4pH/ ��24t3�	C.����g��K�����B�/���.M�Yhz�TiB�Cۀ�r;^uR���^��-�t�2
Z>F�Jz��UT]�2����N��C΍i�}�b����#�o�H �P2#�C�F����t��NQ�h@7A ��6D6�56�m~ w ��X�6��O$�T ��x&g��pFR. 8#���= }T*T�NpNɖ�
	Dz�y�d���\H�B
���`�^v��!~����!�s7f�W	�Q���:���/�H��E���:P �����#4�� ��A�N�N�QQK�1�
�@�F혋���ٌt"������M+^F@&j@@t�&�AA�P�(�ҩ
*�>�j�s8s��ssu�^�k�*����e
T0|�`t��&��_�.<��/���t������&�� �ǀ~��%���Rty��7�1�J>(�����:��N}V��16��
C��"Q��b|�?R�R\*> ?����� ����&�j��Z��"� n^t- J9B-A5M�d|=�~ ���� +����z��
zʇ�~u*�z�����f86R�&̜u?R�� .h5PJ..(���F�$�H�%t	�D#�v��$@v^�x�a {�t݋�~ҋ�p4�ڹ�(��+�{� G�:�,B���� t�J���� qA-�w
-*f�� �uts��l��a&�G�����&�)�^���fW*Z
uS'���.> 	�U8�w��."�c}r4
g���v��7���Z��j�B38F��� L�6N�U����!���"��	!P��R����4����.�[�@��I���*�0�"R0�V�Xa��d���0G
@ �&�oB��ٌ�''-Q�x� ���Y&��/�����&�t6@;��%̗%�w��h�ʀ��P��~.�ی�"w�w���n��b�~�` V$~6�S�=�8�(a�� ������.4�6.���a5�A���Nn�ڑ�=е�%����tb�<��G4g>�P� D��H?d��6��4�r! ʬ��@-��p��;q�=s	
@��0� ��=��tdŶI
�a�@�Q��w��n�
�����u!���&�w����_�fY'L@�#��rQ�5׉s��y7���z`N�PwD��J7@�MP���q@!�$�����z@oy�
T�`�u�WY���%t9�U&
���	)P:w��T�
.Tt?�7�r(��QW���e��������^AZ�Vs����)��)��:
�9v�K+v"�V���{ĸH��t).(P^t]d�E�)��f <�`B�" 4'e�s�줨�6�*"D+F8��� Tt�+�ψ���(Du*\�Q�I��_u!��aQ�Z!R|a�:(��L�v��VHt1
��
��)
w�)��9w"rG�s��)Q�o֐�y��f��b��ˋN�^��S^��R� ����M���ě��w�q���8�   +�+�;N�r
w;v�vȋ�v��FPV,'�
���[[MB��r���I�8A �Z��ʬJ�T��P~N]PFǸ���] )HH�^Y譃ۊ8��/�Vd��^�>�;�;2�k&��;?w�s*1y!wە���b�)0��JJ�V�/�ȬN��L�r�PR��A��W- �>�C�ɐC��1�� �ٱp@��&�H��`2���n����� �C_�B���R�(���QF�V��W���h�,�֙� |ˀp�~ tFC�E��k8	)�Ps([H"�`��Y�o���LF�D	��,�>�T:�#3W t�V��F����:p��@ϗ�����V��R+�nM�@B�'P�d�#h@��,�d���c�,�Mt�P��f�L �N�)N�@/i1�F���]� "�N��� 
�}��
�~Jo��*����ۂ��u�p;��\�IBf�r���⊽t��r �!�$��<M�C_@���	1�'_���иxM���k�RG�-�(F)p����)�LR�|��p�|+2�ҖtL�H�'DID\u=DO�q i(�(�=`"M��AQ�6 8���Q�e
~�k([Zz�``OD�EM%�S�y���K�'Br~��4��d��\���f<2f�� �\�$�x�@J�� �e
z# �u�PP���lC�bQP��Q%X�%�%��R"C��#	�rj:�jq< ���:��V�P�r��V�(:�SpT����2�����H���./�{�#�Yt��h0Q��c�x�e;a����@	�	�A�SW ���9�������{/�|�J�MUtMMiM�
Pkt�qЬ�=�@P�UxP�9�]�� ��� �mD��Rx#&�6���]2RP��Z����&%��[#�P�ts� (_(L�r���/Q�@��� )�&d&�~��&� ���H�� ���+�b�E�=g=�=��R�j�R���m�8u*H����"F����Bq�G��8@p�S@S�6�6��!�sT4{����C�V�I-���-t-�w�-��-�-u-���-��-�-%0
����]t�1��r1�1�z��1��J1[1>J1��1�k�1*U1 1��ހ1��1�1�&+ ���#�7N��T�:�}!p��A
�A�$A�r�"1޵1�*G1
1�4�w1*1MQV��S���JR�A>Z�Ar��r�^1V;M1�1�(1�r��1f1�U911J���1~�g1�1"Q�4z.h8I�R�@(�|v|NK<$I͛��@B@bDfum@��u'�&| ͦozԁHq�F��E-8���� �ڹ�u�@S��gKurX W�U����p~��l�T� ��#Ռ�{L.]]rC���3
�H\�):h-���"{"��mtM�����Q�~�	�\��5�F�<@bXt<u0ßT ���a:@(�L�c�	�X�,�~�Nt!�At MuVx�RXn��`�Vu�A���w�~���,{�P�4�Ό���,��d6	�&$��w
�%�Qӟ,{ G���FPR}�/l�JV��ς�%>|҈H^O-O�0	����!@Tn��zP��/R��4�NA%&�x
&
��d���{������ �uGun�~B �;ɠtӧ�)�~���}����C�f�K�� =��"wi�rl�-v;�e�o<�lc=�K:�}R�]�ܵ�$3��Dz9-P8f8���J�JP�-�t�H^�t�^��HR�R>�jXL�$�E�<�Ƈ��5Lz8Ͷ�m�v^y$ �s�d� �� /����p�����0vJ���)�3Ǆ3��
��	�) f�)*���0),�����%���F��~����B���05�@Z2�]�4�O@6�Ht��E6�9�TH��D� �<t�~�Vu�ER�A�T�<Xu�!����p#`c14����t�j�����<Su�tO
6�u^��B���E�=�ȪPu�� O������Mu$��6f}�#ըNu�JvF�f2��!��M�6$��iA;	ARW��>W�$}z�%���$] �z���X���ju�ί���Cu��
=���Rף�cO��Bb�u���dmʒ.�z������)P��,��Ö,�>ieQ~�p���FsKq��#$R��$u$$�Tw$f$�Q$��4ݖ$zu�$-$��$�$	+�$ $��$���u$$�׵$�$��ݺ�2�2��G2~�l2R�*2]2�]��V9W�$
$��$�u$$�]l��$��$.$ͮ"$$�#�B$���	�v�̌Ht%.7-3��>�
rɤN?=�pz~t8���?���)OO��*P����<�Qȑ
�p��A��F�� �� �P�N��Q�2 ������F�yStB�f��N,�jjP����Q�7 ��/D��GL�u��B����i����$�b�L�&K)Q^�E[;��ڨ���.)s����F��Y�`1b�C�|��M�ϐ�e���^�V\����8�a��M���IK4��K+��9pP�V��T)�c
���. tK	��������DI�mi�i\�vF.�=�&����&����V�Z?Fcr�aO���L R���V�U39Qr	w�	_xow�&�e�0̓� ;&wr/2������O�o뗎���Ԯ%�f.��� ����
0G�PI��^���p��r��Ja�c\��<t�-\�D �:9.�)z&'l���z:>��,Ͼ�����DQ�����JR���w!n�6o� �%���g�M�	HS� E^#�X'+O��? my�bٸ�lƲ$����v��*3S���8��(5���+T�)U����|H� 8-$�h��~lr;�86p1��١��Q��K�F�
/�d �R�.b)��!�;t/�����������f0{'�=K��7��%��Ǒ+�F����~�!%("���\�\	���V�����V��*Y��XJ+��S��U��Rֵ��\��/#L���ź�:dCX�"fm��^�$��|n�n�-��4��Q���+�F^'�6�@��5����ui^P��H��;ԝ�F �ig����u� ���^bl�"�y"�:���|���v�yU{�����e��x�@::�2C���aj����>�a��R�b��M�;r��	 	_ �3�<Ot@ 9�~�Su($��G��IK9LO�,�����(�Gp��t  �� ��	t�i����8�X��� �s9��f��؁�W0�9� �R&�T�? th���-#�"�w  վ��&���Ù���f䢑�9erF p�>�8Htv�o0��sC ��������H$H�^���Vʡɤ"r�ģ� GG&GtJ��P�x�1� &��{�jQ��6�H(�P+�Q��Et~�y�8�.=("=� �jU���v���Hf;B�%UR>�
>>�>>t�&u&��i��>�uUb�+E�+t�<��\��NvȢ�a/\P�*��Eg���	FSq
�ԃ�
�F��h(�� �؋�W^  F= ��	��עt- D�u1�Y�J���Eyss�:�Y$�* .�Gf� ��* 7��7B�����p�'��"d]h,� �-9G
ut �)��!`= t�=
܋�=��=a��=�=�a&�=�=��=!�=$�='a�=*�=.�&�=1�cT�c�X�
Q�#�p�F��I�d��D�2tNu=!C�"�=;�& u'�!�@"��ª7���`N �O��V0�=-b�w,th,	� ,�Mt,
t7 !W���>����u�F���WC4jW'"��J"���"~�r5ߟ��`��F��Hr&p�#�g�$�A��9�
%��3x9�!�:+�3�*���y��x�k[D@(Im)Z_�Yg�����79y�c'�<#~���,���;K,(BO5�`�/��\���H��]��EW�d���%zp� �>�2M� 5aHu��IC8��8G�!C*�����?��.���/�o�����.�J.�U�Q�T��j@�N�)*� �5e� j �a� z���\��$�5����-6�7]���(���v�01�����G@�7��V��(����z�+��m��7^y�7�2��]H]���&������8C�E��<�ƁS����"�=�@+��+��+�A��@�.�|Q��C2�O�x}5�Ex�Dl&J��E*	�ѐO��V��HCC���ad��VW�rJ�hf���Z��J���Bb�J6��t*� �w���.��Z#� ��"�"###(#4#@#��B�tF�X�'��ET6�K�t����%D)L�b���O��$�^�hX��	H�3�R\7҃xD�*�SmpT����iP<���U>Z�၃��U 9�E��;���>h�����nB������x�"
����>644�[��������bt���(��̸cd���@We.0ѢI���)���T���^���h�U���8��V8�8h�l��,�^�j��_�@&��~��(�p����$��t�D��x�\��]�tW!�u'|"�':'���S��F�D)���tB��=/�wm<g�A�2,E2,w]�v&��!�&�#Hr%�Q
"��#,Qn2+2�R�2��,:T*40�	�$\	���;b��-c֒x��@%!t�Ux��鹇H�LR �$Z�st�A6MA�Y�K�pl��ɺ��d��*�K ��.$����+FĐ�F�5{M��
ɯ���Hh�:��!�Iu���%��0�� �!!28��X~����}2�}����<�2-q��iߡ+������v$�,�͵���Б3txEx[��D�q(���S2tA���n�	 �����`V��F�	t���;���;��N���h����ɬ6
�� &�������@�-� )}� p�@7����֞�"��6���uP"K��D�J	N�3R���^K������n��I0x$A��<Ou=��|�Q�	��qI�î����P ����"��A�� #U�$��|O
q%	�,86��?E%����|r ��I�	���۟X���P�ޚg@��Z�)�m��$r�MX�C�S�8��5�������K��A�|��J6q@�3���A�&�����ո���!*�B5�����:�6tp9F�2�Vhz�� Q�A�F�h��u��#ee�"�\F��@��AH��}�0��F
P�6���8@/e�^���j��� ~��v<)Vo�TO���zF	�	t~ü�{3J�9��B�T>�i���
�V��5�^���������݉} v�}�?zPzuϣ�wu�t뱐�t��t@��V�y���ap�E^\ď��: jKG�Ʌo�����}��tNr�H��;N�������lZ�]� �ԣ;�	�����2����t��1)����������*� �x�^&�G�f��� �y���V��v��L�����%@��% xE�0���f^�����yE������r��U}�@&@u?f�%^�������v� $<l]l	7�9)����R��N��,j�tg���p�b4���������������W ���O��+�^Q��W�0��ܓ@$X������uk����PF�G�GtO	�,7�M��w�����ݙ����b\��+N�N�M�}��@;rk�
vM=ڌy��^_!\&�OT t��*���~
 u'��	�`JY�V����@|�H-�"u�~��)�v/"�j��g(�� Z �kKJ��&
�d��O� ؿ�
� V��	=�Kb��8����
S0����  ��� - �� �zI��
��IRa����F�t�� ?��+�N��V&,z/�R9M��s� w
^w4I�^ �^�/?u��:##F�*�$�n�~��EȘ��� ��w��w%u:foq��bWtw.rvGrw&�N a�*�+������&;���Y�G�;��M����S���<�v%�Q���	�.� �,dt@8^b����o����!�a*�@���6�r&S D��!?A"u���^�&^�  w�F����Q���x�B�[���Igr[�'dvZ=�Ў�`�Xyb��5�|z�|��
4͑���뎐����@�\���8@>���ʀ ��?du.uw�L����
 ��� �:��'D����NȈv믺�$k������ � SD����'�&_��p)F��F� �@��<���KV ��@�� V�t'�~� u(�6!W�@@0Tcvh�?u���e��X�-�.LH=�LLۃ~�L�ĂL�	�{Aa t�E0��=��N=Uu�-&@�R�}�F}F� �p��9'u"�,��<�A�.��t)��u��+'��Fj���F�-��h����w���]c �H(=А,�;B{�;0^ؠ+��
�9�c9��\F��Xvꩃ ( � t�두�Ġ&��Z&��� f4*�.8�F80�6P� �Cb2@{V�bQ����SD2D.�W�����J,��J�u4 :4#8` u6\GA�,���*$y@
�����@�v2��S<9��>�te�w�cP�F�Y��hV�  P&�26T' $���~)�N6���'�(8�TL�0�
�����Ե�9�*6w��3)�uT����5F58#�5t�T�P
���(P�-DM�@ �늵nH�G|ή��ô-�O�v!�����čN���P��� ��� /Q!S	 ��OH�uc�$�>`�*���Lk��k�쁞k��F��CT ~v|P Q#�����Ր�T����E�a�?t1�����,��������.Z��Ћ	� �|���%�M*�Pp���F�]e�K�M�(mta�ث�vDU�����Z��{�T�'uh������~� t)Wb�]$3����tt���K�`�%v�B�"X��.E���E�ZV�'	d:9���NFd�DNT݌�f�h�j�H���� =����6�(��ɭ��$�&�K�Hy�6�&����!V"Vi�aO�vPa�띐��{�J�E��u7�Ì ´Ɂ� ь�����<DO����V�N�4R���L�+���\<���c������`_F��k� {�X�{�����g��'�t�� D׫  Rh#�w:�*�
*N���NQ��F/P�(Á�	2�vS����������%����P��� �Թ�ntVթ��P;. ����N�Nk��F�p��:5MH�5?{��56R5�#:5���6M.�6�B�0��2��.0�݌�S���S��(𐀴u�
�׭�lj�]�'e�?������T�/jK�vy�W����x�Z��`����~��up���u�lG	&B:� �Q�����r�40���F��N��򻻪�����%�� ��'�����ꆀս����Ƭ4�| WV�*�ү�  �hk�f�N��<v% v}v��� �8���> �g��~ ��KO4 �U} ^�I^����@ ���F u�V!s�Q"�`�<�
�F���)�%� �d�^�/�Lȇ
���G)����=�) �p�x���� �F�ˡ8z��P�~��& �UWV�*` �!QR�,X�Zщ xF��V�^_]��������.�xmm�2`P��Q�N��Q�-P9�u�J�/c�]�A�c
 �d����9�daqG�
&8t�r�ru��ru��N�\u��\u�	�\	u�
�\
u���'9�v��{##��c&^)&P�J=�W*ʽLLR�&&�.�=A�7{�Q	�:��`'��
�J.>	.0�M`� �n��@	���gٚ�7(�� k��&^BY���%��{˺+_Pv@_��� �uZIZ��s"��� ]�.��@.�t��4�4�94�t&<t�#<�&�eQ 8�>�Nx>� 	+�u~�u�(x��r��4��-W��\��\=�uL�-R��R�3��k��E����)���mns�]����-��&]͈�����&���� Z ��]�,/1��($0))��!�@)���,�,�A�,�������,�����]�MD�C&�p1�nF<PH�J��Ht"��
|�DpP����	
��,	�H�U���D;Ad�� c�5t/W�W�������F�� ��t-B����Ή��=w.O��.�A�A�G�հ�I�R�|r�`7`u(�_�/^� [�M���ع Q���~IY!�^)P��_ �*���ٌt鋪r	�Ur
ɋ�$�u���Z�����~��FQ
u3�2 �J��a��t
��t��s���2��H�P�G0����0�E6��E.4��H��o���u�mS�� ��< �?��/���h�� b�9rL�r 4g�p�G�4Wu2����S�VH����*��4	!QD'���.h�����Z���z��� �],
��L����w6���u����Ί ��F�$�+<t)M�$}��I�L����&�#
=<uuU-*-�$��Du!��$�������� @-�$��#��  m�t	&;Gr�z�SH��}��&�fWV�FR`ծ``�`�F�$rV�i;�s�J[�Mg�F�Ӽ?r���M�`�g@NZ1�@P	[0�a$J3�3 ���0ع2�N#�,Q�����;TO��_� g�]�eEh�@?�5���A*�l$�e�H�U�RM6f�,�Wn�� u����m����t���¼�$r�F�.�t�s	���^�������E~���p �R�����L*���Ug0�����~<u�9F�'Y� ;@�@T��;BI���������;�xtG�  ~��v��Ў�� �U��Y�Ԩ]�b^���!#��%��|mu� 1���]��+�L�N��b����AQ�.S!G~հ��Ъ��������\���T��f 耛o��%��2��1'���S����ތ���s��|��N$�������4�F�$-Q�f��qLiCqQ��[B܃�*0g��L�r������=�`�P^.X�F 9��D�#9GtB&�B�E�� ��� ��/Q�Ը�WU���|�ɞ�@qR�OVw��N��r�������-b�A� ���L�;�t|VW8�7�2b�V��ػ��~W�'3H�[�T"TA�	�JX�ti�S'�F*���FRt�s)��L���VW�����6��;h�t�ȀP>� �S��  �8�ȋ�b�b)��)�4VW�J_b�=t&Bc�P�V�&�� IG&W�,�
�]uӧ-G.׍.
B�j��S�F���,1:R���*�*���^�P�WF�n�*�*d5�eE�Vp	<�>�0uI-7 )^$�7���x�7��܅�w*�q��Yt q\�u��F�)��N��'��me�ԑ�߆K���B��-�:�_����:�E=��۲�.Z�,~�g��Z�4�Z�G
N�} 	�ȹR��_�8	���,�u��|���{��-��3Q��?��$m���~��t�I�������,�<���Vlj&�t�gf��%'
 �(t}P���dK���E��T�cJ���쉶T�	�p��oĸ/-8��Oҟ�Z7 <s��v�Q�^��� X��m��¡l%©�T֚��hQ�Q�X����t*�u�o$R��T*묐*k꜄Y���%��e�@R?Q٨�@*p���<�rn� 8P �9F�t�/~Qэ��b.�RA��s��r�KvG��N� �7v-�>=�u���t���o��q�������Q�V�"`��n��p ����7>��&��ˈ���"T&xrL &�)
1�6"���b.�"r}"@�'t#�F��#�@ � ��X� ��#��~�.�rA���z�r.��Ob
j<�s]���ِ�ʹ%4c^�6 t��
S���7j�jM��j�r:���K#NcD�l�v�-v�+��4Vi7��F>�o�s��x��u!��ƃ�+� �/�0�T��<9<w�p�>
u� �<Ot� �������P�Hp|Tu	H	!��<�^�']â�t(�~(�88�����\̿F��	��v�Gm��^ �$&V^�+�/uՃ�%u*��s�V�L3jՆ�������&����^B�BB,aXWT<�*����u9Rk��P'�o�ȜjX����9��(@�g t1�g* *��
��X�@���7�K�m�F�[���ט�wR5���J덐N�V�M��s�R$S�5շ�W���Ϙ��P.���\죸�d	V��V%�V���d����n���p@��9�1 �����<�<�|%�nu����=�e6 &�2�@�W`�GV ]�\��: ��t�z����U6�x���5�H
.�&ITh��he#KRu�3e#I��u�����dU.�̏�� ��4������{���Nej�)ts鉈����]=h?]�^���\:	%x%T;79��D3��ߒ���>��K ������t��O���� �Y�?H� ��E�H�(�0�8Lt���P�  �����r{��%�%[1�<�x>�[� H��9@.�u������� ��v���U�g��Nt�u�&Q�2
���[�! VdUE[�E�˪F�Ǚ��Ub
����6�������D{HBji��E�'�����V��fLN51��VF�n�t���"��F���� )�.7Z�;�Z_���u�ѷ�v�t(w�"�{����5�W�!��]���u��0mu&���>�Q�����i~��r��a��S����H�81Q�9@M������\ԉ\�&�J�����������m�:�n�9���	 ���7��0��+	0>�Б��  &t%�ۋN=��_x�_�_-���-���፦M� �@�p�I{�O߷�T	\c�Z�>uD�G��9@u(E>��^�e��*p����30� #�A�	��a"���'bh�-<� ̈P�$|��(CF�	�q� 4��i�9�\m�� ���4 �"V��i���m�:���A0��H6
��VA���
� ��/�F��V�4y#Z��P
.
��+� � ����؞�~�3B�B��8�}I�=&e�K��o��ZN8��� �V���l�v��FZ�R�W P�3G���5�Z2r�
�I�x�̈~��չ��٫��D�F� �u'!"�t!tt��L ̿�f��s��sO-� ;s��@@;",�|������9s��}1�!L����*�^�^i�{>p�t�*Z
r�lɈ{�  H&���V
p)��Ԓߊw�dRA��5-W
��� G��F�<���f����@b_�~�Suu12����5Ք����A�3+��vzU�䪖'��'���@Ft�����U-	
�,��xw"!��9��������~"��  P	�D\R�p~n	T�6R���`�
�Z����vy��$E��������StD�~�Ķr�E�d��r��KRN���t���Mt���	�VX�띐$�F<�!t����ƉV�
��Ү�$�O/$�$����� w7�L t
V�RPQ��n� �.�C���C�-�g��]���M�F�*�e���N�֮*�	�W����+�����3#�	��(9��J�O���� ԩ�� ��S�;�ļ�wO��B779��d+҈S�u$�&�ۡ]�E8���)��v�9�!�t��s�)OU�m���z&��p��y��kH�6���wb��~��������N�Q^H']=a��r���`
^'�b ���H"��F�B�@�T����̋:�{���F�VΉG��PJ���w���~p�#�"Y@�u���B��r���[��M��e�O�}����$o&�
����h��v.��Y�M��w��������� t$�9 �$�����L��o��h�`*h�V,hY��ʴ�t$HM
�h�F�E�%��M`�y���(V�q�t�0'��@�����fM� O�� �9d� �yW��� |�@�W�Y�
�����J~'�a��2ޢ2��L��:�sA��n��t�P@��;��;�\z�zD���;����p
$�
�" ؿ� �� v�]��N܄ҋ	!��� ����k�& Q֬I"�$-H�>]s��]��0]��r>ڈ�s��e���M�bR-��B2�tAD��)�v:�]D����^���H���^]r�T4�6ؚ���`�> Ru.�>u"���;�oAw����o ]�����gba@�o�vD�."���?'вu�F��N�wғ?w�B	9s1�yg��� 7PE��*�? t�:��u�<uM"ee0�뙀~*L�C�7���DT���aw�l��V s���D�}h�G�4�&�G&�G�ԙGL�o�L�.LL�Kd_O�
.슒,,����f � 07Z*�F��g]9š������褝I� ��F��
�t�p.u8�m�s2F�F9-vS(�P6�����F����$<t�(Y��l��^g�u�X�룣x�t��wY+]t풣�
� �,I���\�I��G ��f���<��&	����%�A ���% �
�n��+�% TD)�%>>r)EF�)-76��>��\��\��� u�zrH��&��� G����<;�M@�`�� [�%;��!��0��3B�`  u6��uz@��9gv$P�I?</ �U<��t�BT���m��K�"p�WV-�]���ý������^�v0-�� ;&�ۊ���V�
*��H%�$|%�������R��~��.�	2�o;>���Q6�|6��Q����D���o��&���y���I��K�\ξ�O��L
g޿��F� d�� � ��V�C
[S�����9ݘ��]�� ��N�N���#�0�	��+-V�'�30>�;rw;�nv�1#��U�o�P�$t�|���诚 k"��V���i��u,B�}8�AZ�@f�|�� P
�_������f�P<GSw�%�M0q����F�V�C��)�V���Z t�n����_�Tɵ�_F�
F��`!�F�%l@(a�$ѯ�Kt��1R��މ۫�2�͔��P�)�EZ����!�-P��� �̾��+�	
Q��$#V�OV,�Q�NES�S"Sº뫂��f�������%fp��>�΂��9'2)dn����� ����[ %�߶�߇lwGQ }f�.����+Ҋ���Ԋ���=�q又i���  +���Ӂ� @vz+������E��N�����I�H�Fv=�#rh��r�3� �O��0l�F���PRQ�0�p6
r��3�v
=7L�v'�N%Q��J�pw�9�J9�/V�N&�Q-���.�.���-���G0�r&Wt%�%�ɠp3�WsC*��m� Y����T�{��z|[���r)���.�h'�RP%�����L` -w�,���J�"
t��q�p�4\�� �B� t/"��I���Za5�d�����-T6d0EV���� �3�]O�O0�FP�!O�
�*�k5�Ei�I	�s*^-��Q�?9`!�*T�-OMF>��*�6�蘃%S��[lܿC�(� �1����H���B���=LRB� Orwt)N
v;V�"r�
r��dF��9Vr9��[��\+���.�4L�rL�v	a��bGS�6 �6Y[6�����N;�e�t t���1[%RA�sU�����~&����wrq@
s��
��+;_p;X%P�\�FP2]���u$�����.u�`j��` =pIj��K��~	�^=W�W2��j!l��: ���N��+�+�� � 
�t(�����u��v�~�b
 t-�L2%�6N��#F�#��t���du2�G7m�v�se	C]"4$vV��\+�@��ȋ�+����������s�^븓���f-�!`!`��d^4[Z#Z#Z���tư��+Ev@���F �aI@��� ���%�r� �t�p7�u�T���jr.�>�I��!�> �z�>3'5��>Ѽd�
y�U�	�^��^��.7:�:Qn*�,^���7G��|  �vo9oYU�
�a�����+�s�H���t�
�4�>���P�\�X�9*:�O� ��6~��*]���9~VsI� �l��P ��ƃ&�6�W�n兼@�t+O�!0�%�O�n哋 �O�"�xd�l_.W�&��p��:T��s�T��n�W�r�qһ������oVQ�^�i��\�6 '�#F�#V�j̊Lk�v�ocp#&�c눐�=D�u��^�3!���ױ��,Rr��R���V�t+e֦�c&�t�9p�Ю�+�������z#}���t��+7�;\�W}..�7���j7�v�&�?��v܂�J6H�7�\��@W���..B������A��� Wb   �f�!r;a@Q��-�z6!0xr�`t pzpQ
�9�\ø?��=-<������|�P�v��x ��&� u~�J7���~3�T|APEf�+ 
)ō�>}�=u�O�Q�z��{t�9�]������E�
z;�����{ <�$�p�Fw]��#s�0��<�P}#��n���^�T�I�� ��)���"�w��3�}o��=���yL���=�����<&��!��!�9�*��:��4��]�*�A���O ]�Q��\�	+�w/�)Q���E���!� &e6��
���2Md8;��	r]"��J Q�� Rb�b�=M�L�S��SnQ��
�,)�)��  �q�� ����(��� ��Q�=Ttw7- )�t�-�u;$Ɠn%&
PW' �)� �-\>�- ��t�HHtܰ�&J�~I ���� �� &���gJ����
�p{������ %����MI#q)&���WAC�~I\b�>�A�8SD�tq��v�ĉUxw��I_�|"��> t+�
Jv����P�p����!Ɖ�5U�P �NtQ�p5a�w �w�z  �/$o�I7���6=��$��0��*(��ˊSݐݒq{D��if�u+��	�!��`/��@�m�u�d��,�9˃)�]���G���@@H�2K��(?G�Gm�`0&+�84-4Lh-"ǸL'G��Q�!m�V���I�@ ��u�d7HV�5I�u�4wdz�^�� ��=��	*t�̃¬���Ҝ&tF�W
օ�zax.�*�e����F�&9D:�� Gu3�N�f^�S<R:H�B��P�Ҭ�Y�6��^�'��<�^��?Gu'6z�@P)Z�)sU/vO�?v32	�fvR��7<��<�#�\�H���9s:p&�ɐ�;I���Ip�s�-�����������ӌ���G�u�Gw��!r��P�G��VR��D'
�P�G{P�N*�{��*�Ӗ@ ����v�k\N 0�Q�^�i K�U�m�-�X��L��U�d������gt!sN}���1�+p&�X#��*�8���ٌb�[�, �n���mt*�.�t��M������$?�tī\���=gS�!�*�o�c�� tB����&!u^��Q������`<��/;�F;	��7X��#���
� �@<t< u�a�NFf��$!�� �����t*��V�����'\Hc<fR���
(��wc&y�3��Cʂ|��/ �ݐ-� =	  �w���.��	��"	�������t�Y��_*��,	t�u�`��O`ɳ���D�S�~��H��u��p��-��8�/�Z���wl�uPl]�Gl��l$auAsH뢐��lO���$N� 8�uS�^�����?II��(��^#c�t#- �ܹ�p�2+X�@+w��u\{#�	E����*/}�U���QJv�x #�r
�w�n�V���^��BR������� ���C�d�����N#�K����/8�,;�u*Dºt-��%;�VV^L�t!�?��	g���H<�R*�*��?�"2��࠰�-����'�x��!��<�������	�������H�������x<�������������������������x�����<������ǩ����������x<���������y��s����m��g�x��a��[<��U��O���I��C��=����7��1x���+��%�d�N�J���" �- =w v�2� ���@  ��^����v@���F� �Xdjp|��> ��R�КL�� 
"( .4:$���=���� �����v�B���kBF�*��
ݬ�%��"�������~s5�#/Nr��Or �	��;�/�W �N�s��;�q�dR��m�p�@�N��ܧNA�҉�,�^�G�W@%uS���x�@l��AA�
u��ߣ����-[�u��j}`;Z&�Ga��y��K�GE&�GQ-N��gG.R*�-TUVnI�-�_7j�Q*�QP*tmɤ���[t�ۊƨ�V�&Y
��c̣��J�!w��b�+�����6�����V��$g��� �ԃ�&��G�N�-&鐄Ȇ��pqӇ���q�Ǉ�h�N ,*��RP����»R�%D� � s  �<� ! 1wH^�^�u �p_������h9�܁Z�*�S�"y��� d�c6Q��x:]��Tk� k~Z�����@��.m\�@�FX�Ez#��P�`�5$F
����[I���.�w�3�ݷX�V�V
R�����
�4�"������vWV�F@B�  �G�[�? A��rѸRP�[v��tbN
G= u�_Y�0f�+!��'Ѭ��u% �� �vUlT��(�N���@$�2i�
�1ī@%�P�OI����HzN�AA53����C�!�K�ك��`[�w`�ӫA�@�!�
b
� K������	E��Ed
o�	i��-`ܱ+u�@Cא���IQ� �&�_*�a @ޗ�� p���2ڀ�2ӀʀU`v�6W#��fH���9)c ul�2e'R��stI��`�!V`�u9H%u1P'u+*��Q`"	$����O/�he	�%e�w-�bB� �u;Nu�%�GM�M���K�xD�1��Fb�\�YO���O$�~C�� 
�S\�(~�P�U=|t�S与,X��\���N�]8�xV�AU>��	a��D�����NBA�� �iBR/窢/V��/TtEݸbԶ�f?�ZB�z�ZjZ�Z\��Bp���t���L�~�x����+
=+Y�&�MOX�X�	��}�0*�'m=�p�� j���F0�/�C(�5*�Dt�t� �J�	t� *�N�*Ȣ"H�O9y�QB�9���EVMP1�O�l�{�z��� ���µ�<���<6I߀�)b�9\$Fs�1�1�3�D����v3�&w&�P��*6'5���O_�럐���C�Z��V�i�zVV��"8�]�F�J�s|
�Ɛ�B� ��͜�����2Ѐ�2��ռ�:0��+���@05w�DR��Gn�(¦��Z��V@-��Z����^~��2�
�$��HD���s�;ra'1�f�쒪��᪴�v�"�&�}\�"�au����AAA�r
q^��
�����ˆZ�@�
+�y!P�#�Y>��,r(q ��$�OAA$I��e�����s�/]/�0��/�/�M�//a�@>�0�0���@0a0��K0�@0�8�@@*7"��}�U!8�GV��_C���&�\�j���P���hu"#�"� QT]g�x� �Gt>&�w&�t�Rc~!��yt
�wM�8.{Jޭ��eν�<ʂD�,�~������W\��v��H��F�����t��ǐ*%�q����V��4I�$(����DO�!OQ	5�OQV���!CW��"� �X{��S��!Hc��c"�Q�n#:{u�n ��-fjt����{_�DM�Pj�h�s�#��肢�[�(�M"uG0;N��JN���*�� ���z����$
��RC	���F�S�F4F/��F
FF��^
u�V�\[��^���F��+G-3���[�~̄i^2�`��7���;��mR�ip9	:�H2�2���uz^6,�,�C�,�u2��,�N��%�6y=�b�-��t[p�*����Q���O�_M2���
 Wi���-"�rq��j�r��2$2�p�ɀ�N�z$@��$	��u
 Ip�����h4a�9I�$w PM1��¤�:��:����ȴ(nT�t]z?k(��2@2�K+v
�B���
]�o)�'w�ɢG/�#�"�����.�
i#��[���"[v1 8J� �!c��e����<���R*!w�ϡވ����({����NQ���ɥ--�z�-��XR���>�)�^���^AT�H]�@��TF�r� �V��JS�{��@�+G��-�eIA/3LEc �T t1��;��%�ܳ0�;�T�CEu1;u�E���8�
�9�DuH�t.�U!�;{��HN �UDՎWV�_C8�Gs/���P8	�L���%t(��y�G���
�w���P̀~����q����1-h�dp�V
f�ډx�V�;�� R�Ѧ�S�Qח�D��A�]㨸���f
��)�
�� ���#�W�Ƌ�L���n�ǁdG �c���vM�֑�)�_� ��P15'����`�% F��H����F9��<�
��5��f��sVx��;F�w5z�Pp�z�7+tS�
&�g@ q@ [���"��hD�o"� .�.�а������^"&Ġ���h��Q�d(�TA"��I�����H�v4��5�tR$�oQk�Q��RZ�
���D�:]V ��u| NX��*�����i�n
�.s�S��0�A+N
���#�	��H+�
ȉ�x��tU�u�+DH&�d�5L9+L��+7��Uֲ�W�9�w��$�����+G��]�'{���@	�*�F�� ��*�C��R;�8N��AKB
P2�H����^L�V�J�����1z'�2��2� �hW;u�#\;Yu�����&�u.�R�[�l�|�P��R�c��u'|�+
q=R,Y����I;Ȳ�sO��#+����~t<��!�0)��@���^
�B��'��mu�S�aw"���+�V�o �*+��v�n:�r��х]��P���% r8-�&��t!ڞ�*�*}9J,�>w�~,+�w��\��+uD�H��z�{H;~*�W��L��v�O��OhEA.��pS*�T;꓎Fpm\�q
����w�2���~ތF�:I�aގ��M�B@S��N�� F�T�� �T�S�V�~��t,��#�"�4O���@����}%"dP�?���}�_ ~vj��)NOh�KV�y?FF��	t{��Q�;��\I���E�6NN�FH �ĝ$<�t J�y��&� A�L��������ߚ�"����F�_J�BWVA�~���Q@��@��F@�@5�@�#���V}i�4��F栀������� / ��V��~���
��������T��\�%!�@������X��|h���N�F��B�����KS����G�� `���m���^6Rtd
֌�w�ю�kT���w�V�>�,V��!��3:�PBv\�F�9w՗Bf�۟�?ɰW
�6u	*��.��Nu�L�>�D��u4��+�&m�a ��J!�D�d�+'��m��Ǖ��߯'bT>r+�u��V��{�$������s�T��r��KLKLu3��p�vS%S���̋e}�O$�x9BX9s�F�8� n�z��M��m&�&kp�l֐v%�]���ڐ	���d��[#B�}I�3E{ ��
�+�Q��2�����Bs��<\�t�05�Q@�Ѻ;���EtH��
����u�p��\�jHv-n��T�+ �F���#�	E�
a����~����ȃ)�Qx��	(����MR�l$���g8�d#�>ހ~��BO!�oP�
����	B����<�eB��ηx����
��v�����]�����q..5�P�xP�lo �B�p/��Rܤ�F�s+�@H)k� �)��V��t��Y^�� 9|v����Ì�lK�2��K1�+�ݘ���}���%�ˢ�WR^r���3k)L�fI"��t��m8B�����Y���B���ȼ�*!�
�ddD)F2�Y	v9�a������@�
\���?B���LPzB�ɽ�)�=�N��~� u��xl�S t�0D��&�` O˒b ��1��ظ�͸�ud���R��Es�X�a�U�=%�P�)=#�"!��1x
��
�J�&bb���"r4**�8+pێû�S7���Hu,�"�"
{3��^�lȄ_��*9*䨀u= >v���%&H�ɀ�c�7	6��&N�?%�" ^�T���z���F������tU�nz���2�Mwh��ǿ ��U`m�8��;��Ƕ)!�� ��u�u�>t����Q���.=R6�*�s-�/��$��^����1 �/�D�䋇v��x+Ck����d��$���d�%��X�b���(������ˠm��,4e�. �@�:ယ?SuLD� ��/���e��'E�c7E<2�t@%t�	�9�����Nu"zҫV����$�%�0@u��
�~����N�������QQ��A���\���^,3���op����`��(�B��߬m���ê"Z�%��~&[*� ~B�ʪ?Ä��/.�V"�"d�����P&q��s�$p,��X �Z�RP�v��\�����:��^�WVǆ��%.��JPp���R�`�2�V��t����)
'�����H�94�9:�F�����x���	�(�"��"u�-��M �u;N��"(�G +@w����TR��m�eH��] �U"E�M�E
 @�=�,ct���t ���.,g= w'� ���.�������J���Rl�F����(���=x
�w�<ft��<X�{���,,t�,#n��Ѐ�0U;�,u �;�BH��D�������� �3� 
t�|�F�s�^����<����9�=,A�R�P��� 4��. �pT��6$I8��]h�X��=�)Ğ�饲��'g�'y`D��V�.t#�H. *
�,Q*u�t=C1]P���u��2$��@t��E�`�1a���^%5�GF��8OC%Ѐ���$�T�<��1a�ʋ�	l�"�/����^�C0|@�{9~\�?lQ	v�� ��1��n��P��{{D+~(9b% tn709��!���{�- �1 ��N���0u'%<'���;��H�<K��O�J�Ed�;�a�$�@$�y��7EH����<i��],Z�����O�� +8)u��N��� ����p@��ٌ� ��JG�tr�.�aWw�P
���n��1H��s�m�v�&�Gr�=1�d$s�'��>N�?����S3�j�0��V}	�l��� u0�>����	�H��
�N�u���*^�dG�N�v���
u�:�!8; ��
̽td�ƌr��J@:u;�RMt.m�3)� B	u݂ �����m�Ku���??����<����?n� �S	t�����������'�&�MM�G^�7
�jp�r�lWV��	���Z���1^����2K���u~�!��ԘU% ��:�i�,����X���Z:�<B ��Ğ�FI*�PP�Y��!�Y&+��}��M�1eq@e�����[�� \DXWV$��H�af��X���� \��Wǆ
   P�N��~� ~.�*К�=xW�%v9uך�*�=0���F� 4ᥦ{�c�f� ]�Q��Q��\匆�.��0QV���X�O Ğ�w��;� �ƆJ� �7���oI�q;�[��+~�ƃ9�F�� zٌVV"[��&��� 7�F��V��0%�b�@T vg�F�� ��� �t����;�Aǃ�`��A+����Q�a0�g� ~,����F�)F�| � ��p�~��C����U�,�{	qO�B
+x��;N������n�|p���r纔-A�H�顼�,���ι����mԢA��W2t��M+�8�Z�\�E���h�Z��њ,�юQ��D�0D7�,+�9G�(�p�>"* u5�� 87 ��/�+:�FG��OF��+��Lc&�6��^]�]g�F���DV^�͛BU�:��@��.9�LW�)V�F� %�N�-A&��@��7���vN@�d9�1�&$�9D�S##u$��$Iz��x�p�� ��mM\8��8 �n�^�l� �u"�>���&��nV{`��&l'*�Tj�N����ƕ$*$�u!>�)��X�Gt��7�|x���@-X4! �zi�8�"�
��3/<�8��u0�Ah�B@{�S
A�M6��}����"#�~ tO�p"t#%Ic-c�Jc�0��RF��0�+!�!V��FQ�E�h�����P���� ��t&VJ{M��6*����ek *
3��DJ'���$.� �$����&��s������h���d!��u�F��Dٹ9OQ!�ѝ�!t@���;A�qJiF�Q:��"ֱ�L�;�@�dU����&�++?�s��(�l?l�������_�Ej$��暺i
��6i�U u7%T��R	���JFtt
��B55N�Q5"5N�5�A�Q4���@���ފ�>��CA�P_�F��"�2)99p�ȶ2�����B����S97�7"$� :8t	�T5T*�	]���d�Y�8S�E�E) 	�zR*>ug�N� `�SgJ�-�^r-:-���04��
_�
&� �!�v��  �TD�����~� Utwj����x �A� o������������Ե�*�R���RJ`�Ruy	��@P��(NV�1���GAݍC�L��s=�V����� ���� ����h������9޻a}   �ȸ���&��� ;�r
`cw;�v�N��'v'U+�R."݇�^�L -\�+00v0&;Jrw;T>v�ދ\M�_ � �r#w	&���P�r3�%�9�m949�4��H����c���V���v���g������<q�n!	�l=�w l��/(�dt�MA�WC8��L?�?cό4�wb4�sO�ܙ�ʦ$a u��7G�p� ����zHH�&;�� w5r	��G� s,$���VQ��>tyo?L1�닐��	'F�<��� O��@���7��v@������h[)v�BAF�NB�� ?���fB�d�#�9;vY��X��@ @�?u���:-��f�#�g�@I �����~� &t��0���V��F�*�����D���h9ic�9k��69�˫r�M9�r����t���w�d"~&���]��������E�L�<B*+ GN�v�;�r����v�5�5�V3���։F��;n��8���Ch���F�6�
����̮ʢ����1:��'�N� ��e � � ��(V������"H�:4��9��~��=�f��w�~�OS�^09I`���" WV�J�C�� /���MDu���
}2� �I��[�Nn3���	p�OA��|�/�F��S	�??VW�D� �۹7���!_^��r����Ua����!�Gn.���0�;���wWy�ܫ���;��pt�*��w��9�0����-	�G�E�kdb�&�B+�Q`����g@�-�2>z�#��L/$֭Z�&`I0�G[���	{������M�o������-���!-2���"g�	�ٚi�,^���\���uv	�K�n�5�.�&ʙr���	�?&�O��&8��t�L{ G��8u�\�u�\�u�\�u�\�u�\�		u�\�

u�S�o9��qy������p
p�����k��sLG? ��Q���w��r����u�	�.	
��
����.�,,�@��V,��,r�,,��uBB��,,.�]������U�f	 	#�B0$7�l$��&�&�\,','w�))�r+��+-��-n/u�n/2��2B5��7F5���79=u�9=9>�^5>Xi ���~��DIH� � 5 B]��vh���9�ZGI�j\K�.�B]#.��@AQ�N�^=��!�T�Q�ӵ�|\m*뢚z�&��D�
��zI+��R���O��9P+��r���pn�n����S�]�=��6��p�� k����n�n��)K^?�(Α>�zf��C �SɁ� і��%@��&��&�~ t
��Lp�i4�y�!i53\�<� � ��� �I��M lv������(��-��Z�{�d5<�e;gP�j1*�hw)2 ����:���"�"�� 2�t+�&O���� ����+�PQ!WvK��@X$*5��"�G&���̑�~��"T����I�Ћ�I��� @����=OS�O'�I�c) &�w�&)+�H�:H-�)�t��R�^Y�@���/50Cp��%����2@��4 �-�R3 F ���&�>T$x u��Z�
P"8�'�^&��<�����$65�7��;9�9m>����VV+���H+�v*�����x�=��pWV݋e�V���
 �˄`O,2.�L�k�v�+ɉ~��  �HɃ��QW�������T�kB����ɔ +)���F�V�;���ƒ��L�ƉUM�.����Ѻ6ά�t!�}.e^���#@v�~��w��)/�+n/�J4�t3Gқ8�Y�t"3�b�^�~Sa�{��!\F��B�U�� O!]e=������@��Vm(e>nF��d�F
@b��M/>1�$V�t��șT`
�#Ҁ�f��1�����ް��0F}�w�D
T.�$��� �g&ǋ�g���#���	�&�(|���r�* � H��H��we&�   �����(�P�P�����>ZA|�w���}� 5��"<^�~��kh�sD�D��=a�R$�b���d H������>�p/Wd7vA.�xJ+�Qfܤ����Q�{�'fff�hf
�WhQD㯿jNl]��)�{)1z1|�np0� ����NW�t�ma//sP'~���Vr�6t1��ir@��@�
+��88�8��� .����JJ��zS��r=O���CV���a��f�nS��	��E�Dlj^t��������QS��PyuU�SD,��j�s�4��z�m�%]����F�pS���4��G����~���+=��=�.�[�MD�t�r	s	��v�	��!�'n�S��N9jw���  ~� z��;s�6����B:�S��9���=��݋�N�<���7��C��� ���Vg% *������G�&���ˁN$Y� �,*�������������/������iY*��� u��*��l�5�6oA��e�:z`�!��sYNM��"WV�0}2�1�2+��C7 \�� ������\��~�h.���������N�+�SQpxѱ���ȋs�e�Ċ�d��*�D�iK,� 2��^�� ڃ��� SV�����U�\�^���a�N�+�钐'Q��W<���"��%��9DB+�#�Q�KMt3�����F�_�u��ް̓�\I
�s6�~������y�3�D	�	�R�Y	���"���	�@�? t8ժcD���Ɨ^7E�$2$���6��8\���y�%xמ5a�0�(�3~��N�hQ�d�^\-yN�K�q�3t4���O:(��rh�|#�u댐y�4�5�!u ����@[���&�Z �8a���1���|�� g��9�9�6�)�&�)p��3�wdbYT�����1;�3����i����v�Qa�#F�Z�,;>�wn3����
��PRj�]c���,.�@z��T{���c���i��)o�^��/���Ni�*�S�2P��̫��[٦�,A�+���.,m�Y9� ��Ҋ�\V����!��<&��pƱ�F��$ڻG��>`޳�����*g��@
WV���T4+�紅�S�2W�y����3�3�H��1	1V&`�����*�!aП��� NF���3�3��vI�~��''3�%���?B�(f�����H ��$'>!<��L53b�b1Nu!�P�@�@v�0@�܍\Q�4�]�*	롰)�9�u���:A���~0W�qπ rm� Ƹ��^�������(�&�&�+wa���$"� d� �f�]��!d�+�RQ�A���e8!'�PY#�z�(�(��-�i5�,�(ĝ(�@&�3�!.�G6M#�i�@#7rPG����m�upsc�"j���k�N��A�j9"�F�y��lj�Myߵ�L�+�t��i��nh����~
������)�gI��I� ~_�~V��*����l��
�n��j��%=��>O�|n����~&be \5����Sɑ�	8�*����*��5�R�u7���7:���~���K�P�BW�V��F#�r�x�~<n�k ��V0��*�]4�d�^�݈\4tDn{�0�ňD�ab ��KW�t�H8�� �݁���
��.�HB�� �Q%,Ƨ#��b� �N
�^�΋����҄��vO	��pQ!���QZe�����T�6t��CP�� ��9�d��	�y�g��~��-����@1;�u�������3+efa
�޽aZ�#ea��2H��$+��G�&��sSj�R2fR1��/�< ,�6��sx� t&t"�� �tݑ>�  ����+5h�#�`B#}��
��y��pnX�xv��eN�R�@B>c�S��\!0���2ј{��J�b���k�(J^�*렐�Q�֣�=���=��2t���jt	jw	��]Y��X�
:��:�� :D A&����/D/�SH�*�ΡH+;�u;V�B`@� @d:�+�B���te��
T�w�+�v��}^�+�ډ�^=
�wT8��a�jN� ����C��hWVeR�9��D1�� `*����Iۭ��SQ�c϶��V?++��85#�ƿ��e�����C�,tu����y �׼��R�V� ��
�%�:~9�b6ȕ� l�6��� Н�-�D	�� 20��%�ȑ�|� � r�� H&`��r��@�D�� QS�}�w;��:�L����_�0�}
��>��s�H���j5Σì\OB&�����Bdy/��LM*��0�>Q�<t\ 	�v#@t0fQ�T�^�dXP�a�7.a��p]����V1�c	9+�+O��[���{I8��`f ��& }f+���(�(��=$@��T��;�M�� �r���*�DҌ��/ ��U��~um1�	�4P b��'���@"O�@�~�N>;Y���S�����N`<�a�2� �F% =����F	.�]�b�[gF��8ƒ����
�&�#��H�� ��f
jn	�)v911�49����˗��?����@���VG� D�x�)�~i�z��t����]�5U���T�"U�ը��qJ
��#M�j�����ӌ�r]�6������A�ӭJ$k����6Dn5�?1��yO��*X}ޚ;-*
�qw
D�k� �?7���x\Bӊ�V��� 
�����BT��BF�F
<��[�Щ�T�*���f	�� ��� Eg���ߧ�	k+�Z>���3�P�,�%R�<+!���n@���.���F�2�������00���
|2	$�֮��oѝ
aH����H�F��Fu�f�~�>
>c]�>*���)]]��:�� Tf���TgF�T��$T�M�T�6T���T����b�����J��;�9���.��~.���F4���� ����� ;^��=;N�v�Qp)mbR��3+$�-�+����i^�Pi�hu(b
�b���Q�F�b��$b�F5b��`M
M_�E�(P��F�\<}�������@��A	xڗt�I��tɁ#A��� ��}�'$�B!�ل&K�5�3��A�6��g`) ���[����%����'�?����Ȃ����|�6�v�k0�F����~�]襂TswGD�KKl�Y2JJ�8�36���ښ(��M�+�;���u
;�u� U�+��I؜I�o��u^��"�����Yf�Y��m�3"�6B8� v<��#�++@P�|�i�������n22�� ��x�*�0o����=�:*�6��t�@+P�Q!d�*t�N��z~
t)+�E(0���[�����r1��.|��V�3�R�G4++�ʐ������۝�w[����.zQ��J�(�RQw�(L��h&���F���F� � I��ll�_�t$�&�?�� tu���n�1�i<4��gD+$��Vk�y"T�>~\G�)
��}~��2 �
�L��Ś�[���,MA�:uht �3+���_J5�9�+k9�k�\V<�tF�s@Ar��Zv4a zv(&�*���ٌ��uS�6L+J+.���"NN^V�F�������}G`�v�E8��]�]8|j]�]8��]�]]��x]��XM< X}WX��Z�[�I[[܋�Ma�g}G�g��9����,kt�q���)��.�&Q����S�F�A�j� ?+`�P�~� t����*�*H*�^��r��I@-��7�;(sѺ�r��$��Ё	�� v?ҁ&�^N�D�Q_�_Ŏ	�F�P0�k��	��$<u�?�K_%�� �Щ���O�GR�*{�IPXN]>n��
���B坾RX~U'XXu�BRQ+�Њ~\������
S�w:�JFH+��'��i�r@�
�.��1�$u��Tʴ}�I�M`-̸�����!K.y�N�8��L�XXO\h:��7#��rnjtЁkP���
���Z���^P֒�Y�l��1`�`��}`m��&EnW�5"�<��K�����vQ/�����B8�F!�����
���f �)�-�2Gh<��) 2�� = s
�u��T$��'b|��Z���s�`1�e&��ϣ�	uE/_��/�/@����.���2(�p>:��L):� w�f�bm�r�rr>p>t�t"���	
��/�*uc.�
�G�d}ښe�"�nd� Z���LR����@��^�����?I�r9�.|ʂ��rE��K�9Av�/9��ЎI>�"�^ت"�
QL`�ij	v��v�s6�Ᵹ�s�
�`�� *5���(����w/kt�:>���G� ��濣� �Þ �><SV7XL��/i�f+�X�-��g�	�5�ËV=�9�8�8.$[xu�k��Te�r�q��U�� ��4�m�d"d
�W�֌V��~��
u%�r#Q*�n�傧G�2s��
 �H����o$�N�*q��ܘCUN|ц Epp�����<�^����t
dH�F���v� -�w�^|X8?��N��mq��O���%B�:��L BZ�Z�3�?�4q��y/�.�'9w���F�w�k��,=�0�
�s��R��8:@NQ�skv9�k`��/�^r��$Q�CIN
QE��� 2�[�o66St�r��. �ގp ޔ4Wr2�֜���,^����Z�1�����3����o��_�F�P  � �Q�y�z튽�&AlV��k}Vȉ.(�{��A~.jdl�l�)�P�"�������U��7�/TڄfT�6R�N�T�k�#L�Z�$Z�O-�Z� 7z�>`*B#��Af^t�aZa�P���IC34��F��;]t��.�$Ls�吢Uj�^��.tb����ɠ`+S
	B��H�Ӛ<q�*$���Q���Br��@��v3��3�O���Of$?+*���b� �츇@��z]�(���FTN���Ԝ�F
�����|�e��b�����j����!�;�it02n6&�h���V��a�eh �����3�{�U!�&��r3�P%A_% K%�+��jT��
5���%�خGZX�>H�j��z�t16�e��� �e��e���N��A�Z����I?� A?7�h=Pt��uB���$����"�RE8����z�@����	���f���	v �+F�F=`$�.���:�Fht�V�|t���d��FB}��g��_^ ��N���Et u�@3���AI�7�,�(7F��l��H2kÖQC e��L����|�%�.�<|�'n< j)���xN/@@�ٙ+�����+).�@>��%��Q- ��P�aVI
���vV�F���� G-(X&4��K
�� � �II��<22m����IB���I B��.�����f @CIt��)�������. P5�Ǿ��p��^��������t@(��Xt�n�H�D�+���Й�}�X@�Xt��X?�td�������
�H
$�VS�^� _�p�v i
��	�����)�!7���
�
���
�
�Mn
�
�
�r�
�
�
���
�
�
��&
�
�
�7�
�
�
��M
�
�
��%
�v  �= w'���.��B�� ������� �� 
(��Xj<�v����HtS$! L�E�(Z��FnnS鐂\���0��u���Đ	�����V�ᚾ~=|� ~$$#�R� @�0�������NC�e�0*���gu�R���-���R�u����מ/��|V|fF�	�$�����0��ȝ/RQ�7�'!��z�L�!QG*�S��&�ҢOH���SB\��ǔ�'(9ŸH���K�ԣG^ ��CJD�P��͈F�<MSBm�W���C	B<�G�-s�C�CtD8 �>!� t>R��gJP1+��{�#�#�@�� ��4�� 轌 �U΀ <���G�e�~��1'�.�M�0�rK~U��PEOG�nj�^�n�C$oE��<���R�t���Tƒ��&@����ǌhV����x1�8:s4t��(�65���ˊ&�d@�-��@��������9�'hO� b��9
LŐ�� ��Q'��
]�ߕ�*D(DW�)��P(��q�V��z�_����lu�ٞP��u��ř�xht�#Du?�����A�p�ކ�-�Jm�]oLp���h��Fu��4E���6 ��G.f ��uh_��4�4m`J�n��fu�T���"y�k׾ykf�B߷�<XGR�Y���5r��i��VR�)�E���SrǊ����H�,7ꬎٚZ�Ш��њ�d�u���ՙ�
�ye��D��g���ځۚ��C ���0�^��&�P$BQ"������N��`��Q��&�A��S`����S&S@���)`�����&84� O:,�,���	&��)���=�� t^��C�j�F�ؗ*������yJ%8�@��O�\?;:u�^D^2T^z�R�VC��,#�0z�e=2���̀�Fu��#Dm�Y(s�^xQ%T���|pQ���~�.X�w����>l+��7?����}�I_�կ�R������Tٗ ��T�����%-���XI��b@��# �$,��*�Z��vup��c �`� �4�$L�f�%�"L}d�e-���a�Cu�
b� �A�l:x��]��-�Vc��c�?�@d2&3,����[9&Tp�D���c c���4u0ll�t9� ��>��S��}�:�/4�v{:�x�tW��9�$v��J;����u�PB�i^O!BN�-Q�
>���
V
I�bK���f���+C@�M[�@�Ji��Qm�F7���� �REKe�E�4�hT�L]h�X����+�^Sٓ����}-�%,zV�Tj��T8C��h������Ȋj|YLPJ^}�}TU$~\2XUWRvDU�E���
�d�����	����:�_y���� ���g:�R�����QRM`�Sڴ� �L�%����Q��
Y=H7[o��[ z	���\���MB$V�t:FVWR� �U���L��	w���	Pr�p9Q �	�g_ ��4�y�&��0���W�NQH�HȩTغ���`Z�������~ ��t�BW�LHgRP�I.<LX<P�Sxz��ED���QJ�v�8�]��vq�1-�EHB�Br%pX�V&�0X�T:���9��邀꠨��:�TҠ��XBj�.�dCȸ ���N&� �Ě����^�D<˦�~=�,Y���	��ZR����D�>ʛ����S� Ɨ�OƓ�و�*u��p�
����FԈ���ꪵH�D�]���Y��wҳ��e�S���$�
�c D���g�3��""�c�>xt!�&�.% ����  u�I"��������[e�W���1N"�XY�2��K����m����7P.�GUW�W(�SWWt�׿AVܑ�h�T�b��;X �>Í�@U>��T�FD�/�}*+:Ƃi?)�u��"	����C�PoQ/�T�
d��/���"���4茔Ƹ���LG�-��6u$�-Q��N���$.�RX14Zs�� I�#Dc�ꈰ�Q�pZ�x�	�CRh�Ev	���*F�z~�)X;Sn8Q��8���T�BPhK���EN��Lz���4�%5烢�[��V_���F�f��Z��B[=/e�2��4�4�KU4[4���4"DQƸ�;�������Z���\ C�ϐC岸���WR��e�,!�F�@��F�fa��\��P�H�E�� e�����L�fSuC�S���� �Iu�� Yf��o��Dp��i^��M���-r$��9�W�����u��~�)�vtpL!9,�p�q����) �	�Fo���lo�W�·���ʖIo�tZ]?�[N���:;���>4����@t��KZG8�B��z�SLLh��F�B:Pr )�S2�����@�`%T$7{�T�W��hOJ���V/ϬTa�c�V��o7���	P����aw"��	]���wFm�K�%-ƃ��*��@u'��b=2ߵ=W��*��Joa�T�&�H	H-�O(�(iu��"*Ї�rV��QGu�s�� H<t�-<Xu"fP8�B�@�S�"�q��Td:<:������R�P5�%��8h����;H�*�+����C�:� ^�@�:�C��0�~
�S�` 5�;F�5&���+Ky�U�#I# �_�0Ҏ�	���<CѤa���뒆�x)�LN�J�L�Q �;�}i:�����N ^Q���R-N�^X�n -W����� Z�w��6J��i�L��[Lvn�f�U�jU�	;!�	Z�4B	�Gh�Mʠt����o�cU(j��(n5�r^-e�rA�c�	(,�*(fR�E"o�h��n�i}��d�Ҡ�Dݒ��h}��3���"��^
�uu!C"E܀\r֒�`A��!�S#r�U#f#�� �*�xR�6Vs-��ڨ��D{ĊF� �Y�~ t	�Hr$lN	��N��tՖP�ȀU��RumȄȕG#�ۊ�W_"�l�2&_�,���x\�u �� q�� �@
�U
�q>}pFF��pf��qfR��(+�$�$��$��$�$ A$��iؔ-ԐD�*J��ot�hx 8�E{aTs��qAw���qN�-'�-��a�s��ND�b����H����t+&w���a!�s'�㴘�F*��V��,�Y'�NB���X��w�V�׈ZD����+]�E�p�}�\���ӏ�f���6��B2��<CtVP�rd� �]�D��m2P����@.�� &������Ċ�M��H�~�~�իa���� ������ُI3Y�>��.d�t� �Ϣ�u-�(k_ֱ*1�Km����':�t�^	��j�*�c�c0~��u��:muk#:�uAu��#��O�ιܰQ����~�tS0��/!���Z&��5d�\^������(�檀�j��nQȽG�
��Q���br~#ve�Dh!��}��z�Ht}:6���� �/�K���P Mut�w�wX}��B"&]����(��tq��  WV�~��-�Ў�� �] �M��ª	.�.�M�~�u$Ъ���&�Z�$w�j�m5E'�DJ8�Q�N�QZ��b�kiF^�_4V�eT,�J�UIo�o����V��~@��n����8X���m2�q����z�z�������}��������x����d��Yu3^_)ώ��F�8$��V��ŕ�9�Z $=, t0 w�,,	t#����^��0&�q��W�RP�Jj �Ŀ�Ȑ$�{��!�!��CC����,���2�X�o�s-f���TI���$�:�oPo	�\���F�v0^���4�t"���!�V
�n�a�ܤ�	�~��kL'���L� �$��Z��F��P�6 ��D(�o�~�5x �L���n�p�p�f�/�}V�t�9�=�9p���l����WV���� U�J�  �/�����=��u � �.� s]^_�6T����u	��Ӑ�$���^&�U}@�urつE~!$����
���o�{) g{���t �yU-��-�$ b6V ���-A<��MO���
���
�w9����S����A�&�]����PJ�F���@1�
�t!�"H�FuJ<�,|^��\It7T9pb�ʉṼ@���&�G `�zw�!�[IfL�����&9&p�͵&o�60��zQW%zXzQ�*=Ut%+P��,*,<��,|�&���p�� �fu�QW14&4^8W�&V@
|�"� ���I�uT3���|�~����� ������l11;�O
u� ?���0 &��������>�>�� +��i	� ������u�� KH��^�ȳ���@u`;V��v���x�+�&+�X�#�wj!	"P�?��6A��_�� k��
4+������9�f�)F����������B�evD��^D��H? =Mt��~�r� D'� @-���38;6s�늤2�9Е� 4��=�"+�-��R�PE	��	�v�9(���'�0���� H��$�&��C�����#�� QS����M����\�SD �,ҹ ��=	,NԆ���5���+�-����t�l�t�o��B( g`?��~� �ri1��r�B+=��t���;T��W	�8�8v�������u��C1S٭c�N8>� u\�&���)�Ɵ�ƕH�� .d)B3t��Z�8�C.45u�vr@�.Dp+.5�ʻ2.�[$�_�V��A�e!��KYu�}�`�5���VO�!�I���k""�x*1;Hb �J q�������0�W9%KL&��*N���T��}Г�t��8}�r"�}v-��xO@w7��u��ΐ�v'뱐I=R���ߕ 7;)�u
�D�.�b�� )м�@ �$��	I_ �% �/1�*&���)t r7�������!+�L�L�7{8K.�I���&p�>��ptIJ �5ӠG������@9�Stn�����i %�,Ԁ"�W"�V  wc��0h������ ;@��F�P��5���5t`@��)�:���Z�ZO2O�a<t�$�Z *�}�H�eC7�$	2� i��uG�F�*�YrVV_e�9rpCט*D,�NM��!$&�À`֍��^8 ��,� ���=��>=t*&��(�,r	F*An �;vo#D8�R��������,aF"�j���Ff��>IQ�>w��< ]��f-
�:^#)�����?�9��ԏ����
�1 F]V��RD,	
[���؋UG���2C[�W0�� �ު@-.t�&�Gu����bYJ 
ճ\\d^�f�F��f�K�
�Jf;� �@ٞ�F"? "�z��" �3ML�p�v)�w}L�c�Xj.��2�I-A���>(�r8ms���r�a����0��t`9qhu�����V�&�q�$4ɀ�P�����N�@RA$��8M�9!!�wz�2an� F;�vd��&+6��B59�B9�N
&�H���.z1##�z�##�����#6#�A�&� ��uȀ���r�tN�r� � �r����O�|�U=f���0��A@�
�v��;�$ES�^��˪�����܊����B2��WV�T�r0�6'��� �"~��|�Cz�ȋ��z��*.p�c
2K7��	SH ���~�^I��F��:V�.I-x� ��O0O�S�O�OuMHA2B"����)�*�K����f��t`�;F�wB�%����	v�[���B���r3.9���tn{��R�:�r�IP�J�~q�p~e	~W��VRS�XB�B�H�N�V��P�6Q�>  ����� ;�r
w;΀Pv�׋ΉNI�^+�}��b+��l$w��-RQh�k���3���@�����!9w�	7b�Qq�y���S�����u�3�T<QqR8����8�6��0	%�2	���F����V�p�>+>�s�4��$���}�_F"��K3K��<A8����'�:�Y� �U����6Q{�D�H�ſ9rcw�']�	Z��S���EU��q��ȃ� ݌ hڜ� S ��cZ��������uVV��(5��,�\uR�HH( ()t�2p6,8��&4[s���D�~��uE�ɈF)� �|��:d`Bg�6���g ]��8Ld ���d��+4�N��D� �
�À~!��|��B#SJ:P2Bܪ�N�O��+������VQ �������a(�a*� 2�����	���	� "�1� �Z�1�Q!$��=DSu�}!:�T�R�$�ui�D � �N�Q��
 K 	
&����0V{��Y'BI�B���|B��n<H�b �o�����F�T��;��G7��S(~�����=�ɃC+0]����������l�>��*	GC�*[HSQ���m�\s4=����F0�͚�)��t�:�O�*�^*�0u6p�{�p ��� �o}���H�� {@a%lt�@"L=;Ɩ2Z����% ��5��Ӣw���ԧ+�SB�)���pV+��Fꉃ�釟@ �B]l�F�5�\9��j�pg_C�#�<6 ���c�u`�^��Y�W����B��R�>���%9����T��B�\���E��&z�D[b}�LuXa�**$ �����/Ș���K�E�K��b$�}�/�	KUBJK0�t.]J�7�rw90LF�v	�!@~�#�f+6�6�6�܍�> �tf&��aF��$�  &���� ;�wr;�)w-��9?���B:��vj5�n���Bvi��G2�[���r��#>�R�tF7�DpF�+`�p]w�r;gw�n��^��r>�2F]��>/]2�.���eO��N���5�z���xG�ca
�
 �1��C�[� tyOp�i�d ���v�6��R2��s�ܜ����~y%�/�(UI��r��;; X�F�~�s��[=^C�XV��*#��(�@�*��u��I�
�����iđG��Ʒ�ƣd�Z���^�e���a�a=M��&����rԲ̾������Eow��C �@us�f���ȫ�?��d v�H	�4�������-�<8���2��#;u����G�v��~u�H..�� �!Ru�4����S��^-�LV��!��s[\A�p#��4���O]� �@k�R�8W2��*ܲ6� ��ݪ5��uΧDu���*%�$ 7�L#0$� ��sR�)�T7T<pBx�� ߠ99$*1�K7$�$D�QHtK� ��	��'/u6����z�x�c"�9$�v"�P�5_���uT����	�ژA���j��I���념l������V�Z8u#��x�t��%C���1c��
ud�f�l)��~| t�O�$� ڙ=��s�'��Q+=�t����2���q�ݤ:�����r��,ty��-C�Lt@�LL0U�?OԦ0.0��*!��
�%u��C���z@�z<�to�v)�����b�Ģ���+X
/+t�g�a����F�6a������#�f
����&�$�,����
��Hx��p��	N���H������E�,=�m�۸�)��u��o���z�AAv�� ߦj��۬ �^
?#�И�،���D�!ڌ�&��~v��M��hiT�����^!�!�:�2u��{;;��9����� �L�'^��F�9mu1�7��M?� >6v  � *�Ht�H|�H~�H�~J�Z�Z��ؐ�u=�I�tv{��q�8/�3Cf�#GT��PW�LM�A�]R)R�tR�\	=H�^�T��
���ev@ȓ�M�D�jV��. �u������m�$?�u?ߎ�a� �� ��!c�+��jʭ�Kt�·�T.�1�R$ ��R*�~VU��אH������7��D&�-H$(|�!�#��������"b�2�@���<��K
s���Z���L�� sF	t��(���j&\-��>�B9"��������̸^���m�@��`�c�O�j	�)�u�!��+��3��g$������*��	*�ؚ~�����{N�wU�{�rЮ&Yl<{I����F�t͋�~.t�]�g�iŢ�P0���>aV�EH%��.KJ
B�>�_����i���d�4�u'��'���@2H}`�H~@�T��#��r�`.W�r��� ��F�  ���H%�q��O�:;5�+�G~�v�KPN)Tsx�Q6p�����Ёކާ/,��(k�T8���W��v��M��t5�w�M�ѫ����7�؀!5���^�R�&�����Y��&WV򈌱��i�����s�!��$N��i,}�,���\s�^HJf��$!��B �8}���Ӹ���M��qBM�0$��݄�LM0-V�J���t���,vG��+ 86N�'6$H��"���:Ppn"6rc��%d���,�
 
*��_��Z���s"���P�L�!@5���1����eP�zn��N&�{�R�|R~��6C����,�ޚ��� t4��S*�Oz�f>z��*4_�,n�2� Q5Q%R%��(�Q��jg07�2&�G*�=�VrR��N�-:�-J��=�^w\$,s��8����&plܡ�B�[v�2Ө��P�@ ���LP�Lrwݸ4�����K
�(w㶀��`N��;ʑ���<2��=22�	����0���ݽMf�JM5MM���.Q�jN�.RQ۱Q҃U{�� .��O�:���hzh�F���t<�xTk"JJ��PF �F
)�^L �u�R���P~`�����4b�;S� bHQ�H� ��oH�uH�H�j� HH)�H�H�?-H�P�:BHWQH�H��� 2�
E����HHGҟ�I2N�����p
����؉^ ���F*�� &kf�k�1gk�;�k�Ht	���&�R�Q?<�oVS�Ы�Hu9S��V�4RR��Q�<�4�� 
� ��
t@h�ll6HH�!I�^�dj�dF -=��/6���6Np��.K�VY��6��%�q�S�hO��o[p��1�D� ��� �T�z�u���&�6��=�D
���� N� N�Ht3��ƹT����
�����{�BB�cx�s���_;�&.w��V��yA5P�`	)�A�-܊^�*�SH�{�,�/�ϸ���xp�P�p{����{�ظh�t qj��烷~��� ������PJK �< ��g�K��쭸d��j2pB�&{�-�Ҋ���i�F��L	~�]j��HNJ��J��җO@��@I � �o�Ժ����;v1+tuk���9r-+Je� @ J��+�KT�+t�3�	�v�Z	蒖	�	|	�~��t5:�}����\A=��u~��
~�~�3�Wǐ�&���)r��Q��Q_��szt�~?|�; �Ku)� /iv�/��z�n_���C��� �9:I�u<�0�`>}���F�F�[�丩�� =�������X;��P�sɳ�����Kf�	�=d���.�[C� W����p�Cs��f����5�q�ѧ͒��wY��u��mC��^%�S�6O*�������,* ���X�NUQ�n�����B���@m�}-�K�vX�rEJ⦹<���u'9NDBz�/�K�7e��]Q��C뻐�'s�~
u�/�� �R�!�!��Pz6Hu.
JVQD!�!�x��(R��U�b.r�
 �T� B6.��k�8E�a�$�'(M�� ��"�q&���''u�D�</�/qn/���઀��L�7�T����<jU��5�$��������&�T~�T.�E^V0׋t,�	�7��t"=���L��؃��$�p�(�p�� p�5/���
@J� s��^9��#���QM��)�7$l��l���>A"*�ACA���A+x��*]�**�4�*2*��@��8&(��L�Y]B�
��

M
Ht3�����+��l1�q��/�o%o�\wꐋ����
:"�b� �J�  � `Cu��MDu��r�D
v!�q�623�!��- u	�o��(3R�0(��*ZrwE}=r8 �8�D�E�S�Q@+$O+<R=''&WVD(��F�Ht�K3ێË��5^_�9��> �
r��*�2@� 5�u(�
�
>V������A����t3���*��� ���7�^:�$�F쁳ˌV��Щ��L�6�D����`�  ��D�^�C�
 � �V��^��!r�~��V�L�(�H~ª<����2�� �//~��o�=crT��.{9/P,Q�|*�t�o  ���r	��鬬��)�@�s�d(�V���| z�X���*"ø&�&��y!�������tv�Ă�(�S�z �)�R�S���k8^��	 p��VǆV�߳+)*�ݾZ��ĞX��x���Z��O-
^�`�D�PR�-� +ɋ�� ;cK�v�� $T�Ht��þt����9��&2���(�f+.�P.�G�b��6�W0��v�Ƃ >Q9�<<�Su�҃n<~�O9vg���sz���P�����-�Gx]�@���`�y�B,rn�^����\/lR;G
����A�Jv��øM`벐�N/�즧O�<P)��fS�|'$V�WȰ/�W�jB�Y�\}�i0"_Q��b�h{�F�@�73Dc"hړY��g8�^��w�if��n��-5�q7�L	���4Wv2��y���I=���m�O��o��{m�Ruz�5�|:�:����T�������7��u������y�s�FB�O�f.�#ff&�M�Gf�A�;�-   =. wf���.���� x���"(�x.@LRp<�����<��
$��X^rx���������!����\�TPI��0��n.V��`��h#��z��&�	��$5�����������2�� �P��4��h�����Lu��BS=s���c �-��t@��41�	��G�:�����K�N�1�
�v� ��WZ&s1�#��ƟR�{ې����6g�-������&LKm^t1�.G3����ɜ� �y��H=0 wjx�������r�Ҩ�Ԕ��ʨ�.�y@�̪3o���{��fl]�fl��:K&f�� ��V�F�\I��2��� ����d!�B+%J<&���z��������V
�
I\��O^�f
trĞ_��=����rP�o�9�CR��R?�*fZ��F�AG��&�@\'�h[E��V1��t��U��SbD�i��K�D8Ek����ҽ�G��Ӭk�>�#9:��v�b��!��o�tw�l]6^V��Z}�bT�@"�*@�@�*@n��.��.��f..�Ef�f	8���8Tk8	f��.�.&�O���@V>�F*@G��_@��Ё�0��L���U�n��\.V�W�z�;Ft�D;Nu	�nV��*C2�� �4����v0B�ޢ�^L��F n�.�w��*,��
zz @nn* ��no�5�����An�tb�^�/�n��n��>�n/_(�yCC�v�i����+��,��2H�{�&����#��2�u����H�uNJə/���-icGo��@���m��:pX�/p��HN�]����_�y!*V��0-��S����b��E$�\��h
C�vۀ��D ��w ϭ�..`�v.��.��.�Z.FE�<<$<��r<< �~u��*�uQ�v"9�B��Bz}Q��}(��Q�6�6D��6c@���T�?m?�h!��8Vqe��B�-���������� H�5<���P����(���U����� � ^>���r �q���	�� 6�j"J�/B/��}j"���#6��6��Z(e#F%��.��.v��d%�,:MT��&?��?7m&vQ�(/p��/z/(.����)J�888��U8)�+T�.
.��W�+	AF�,j*���jY�_�,#�0�-���R����U��-./DK .}׼./BL�608���]8�803y8���-W�-	�&*p�F�7WV�>�/����
$
q ���/�^�~�9�\����X��ع	 � ������ZF��`�s(P �-���@!\��2x�x)+�") )iJg��  �[����1^3O�`��tM?��QðH�b�h���R), /��e�^��}E
E�Y/�G
��gQRGP	R"	 	 W�	&�	����4 0K�Z���[�n���V�6WU�$��~��]_^&$�� i��B�B���b|A%��#��_]��^J�Gw.��&v�!��u�����>]�� �@�.�4`T_`��#�uT,�M����ht�Vb�hU�\P�UD8v����) H= v���u �������(�2����@ .�>�5#?/ ����x�$�<�� D��b�  �� ��^�]�t}~�*a�]�NBN��k�l�����������@y �� I.w��c��JU�A��&4W�'�iM�)���F�!P�|����")@�g���('�f��໋?�z�k�
�`�]:D!��q00"«�Wt�z#-�P��03F�/�"�f"  ��OO
@���\U77]���C&�N�3��2HT%�>�j.&�3
�v�|
����8�������Va�
�\� ��~��n-N*v'V���?Ad��E8G��O P��V�M �5 �P�f�����*�9�KdR�� ^If�"�2�"����Vߴ�	:/ҋF�̈́�*&:	s�O��h��'�P �{��ߊߺϋ��ٗ�]4��1f1��ȫ1�
�t���mC
P��3
NGP	::�
+:
+2
��P JH��,ȴz�%�%���y���̸�Y�|��H�]�H/�b�D'�D�P��&��s���qce�������V
����{Q��� �RQ�Q�N�%�~�e�>O�͊~~*������m|�v�;�c	2u�L�k��T+m� 2�$h�	�	 ���2��S�,�~���{�z�U �!�v� ������ �i�^����O��d�.��0L��!���٢  tH��� �^�@/Z �x�9r�c#�t(�W �F N�88N�N�i��NtN�F)�&I�]<OO��G��.�7.��H+=�tEE� V�'�MZ$HO.-
X
��sZ� ��^�V��u5a�*_zA�-����
�+��;x����/����!��&�qN� ~[�<@	]D�� ��u �RN���SS�%S S��
 	[|�	s&� ��N�hA�� �FFj,4���#Aj�<�j��"��Q�P��	k8��Z�6§�l9�d
��_�Pe�PJ� �%���V���X�26$k&U�PC�}��,n� 8-�����v��@�����O��st��j^�=M% @l(�����L/e`
W�ÝMԆ<Ú��!�z� ����e�eQ+�R�e�f��CSB5f���SfG����"S�*� {��c�F> V�\N�ʸ�:�1�!���ZA�A �U��/ ��� ��,��k!m( �u|$썞����i�6i��1P%^(��d y� Av��q����^�K��*�� J�o�6���&?���BX�J��S�1I����/���@uD�>�D�"u���*Q��)*���� ��Q|
�2$�VT�˨]3Z�W�Z�UH���o�!+)!C$va�-�1� |�`1+'e<��|����L�V�I����bnD/�:.<H<T4�����9�"Vs~�lʹ��b�(�6ޚ���u,�� uA�$��?UNu�DOu1� ODu		� N�Utl4��F��%]�H+Ah�@��/D�B2�*���$&�w�S�E���=�=F�����g����1��+�����/T!�H'��]�
����6w��M `�&�o��-n-9��p5u��*s�Êx�\��P��u�DJs	¡���v�%v9��29���Tz (t��?vZ�-*�c�<t c��cU �6�pc�A��z�!|��kU�3��� �ރP!!- �ڰ���9j639Gti�;S��H�ͦ��\W��^�沀e>Hut&o��v�d1�r���n5���:��z
�a�(�0��ybp�@�� ��K" ��" �T"�k�]�d��d�$�tI+�S� q�Ux�)@R���# ��v��n!  ����� wPrQ	� ��sE�XI�˸�����r#�P�ܿ�ض,6B ��a�1��+�Q��P��R���L�*e0��e�HT׸�r��xr�~� �Ut�E]��4pLmh
Capx�\�g]$%Qe��]s%7<t �)  �~�Cu"�{�������V�f�3�p��`y�r��ː!5��`�I����u0������t~a��F�B�� ��%�x~���F� ���$v�%%t�{�%��ڬ�dB_vc1x_<lZ��m3�l�u
u
		�f����a���8x8!�v$D�%C��UD*�f��8��+[Wj0-Q��-�@-N�>`  )%��I�����!	ʨ�V��cN��>�v�����#(��-��jTRb �0�Q	��.�3f���VS=�S�`�jE����J�Fl�7��/:��ؠآB)�� �(Y�Y��Y
�ʴ&K�la���̤<Mt�����FxФAt(TBt"�/��$2�Ő.u�"d�����:��I��J� 8���Cn�WV�0 ��UN�DO�F�OCD�NU�&[��B1�.x�ñ��� �؈��)� ���	&����&��* �,tK��2����V1	�Vc
>��� ����Y�� 2��F����|�3�h@�ӂ�������"��626�Ŀ^#%RЏ�u,0���V�9B���>��Ϯg+�¬�..K������*͓(��E�ϒ1�0��X�\��ڢ$��P��o�/�局���T-��h��~�tq��*-�P
�«]Ta<��� id�!����z�V���yWh���	!&_X}j����v��i�0+�y�.�k��_����A"d�qD�^B>� �R�*������t���S���Ū��J�V��J�;�W|b�"6�����a���6�F�b�����̉���L.	���������T�	G��s*�v���z��*���*2�=#9,�$��� �<��it�"V��i��i�	��� 
��`�D�HD_��խ�Z��h����� �F�<Ct@o��/��\�7wn��*!��*v����݇*�"���N��u�FAB�Y��� mKY�U������w_�Q4w����F�F�� �i�_0I�7�����0-I�EM�c"E� 2�v�x�;�u �\;V�uW��x 69�u3�~�u-���V�95wr �9Av���V� 3��������@�f����!�+A�+A�=�0m�AW�����N��1@�t��AA���Q�6d�����I��@c� � �b�:)�Jt�!�a�}�Hg���[2Y\D|2��K��/0�	�@�ь �'6���W�0���`�ʤ *B�R�N�QJ.Մ �=��8` u+2u��Pd\f��*��^7���kk�HR��%2�돕��t#� Qu;Vt!�!�"�~
�z� ��}���e���`���u�ހ?u�}
��9Τ�*r�=���N�H(9I?t�uО[ӡ������(żu��r�ߡPX��u���J�~3gJV�{5�W�vX �JѧW/ȅ���~T , o���
g�$+$�<juZ*�@H�N���������U�V�V�)�����c�; d�
�t���
�t�dS�d;�>; U���	 �
�Fϑ�H�� �$��Y�d�� �1�
��)
�9�{�a��~	^���܉Pq�P����
u f����
S����V��/�'ސ����8W��d�\ ��T2tNA�@�N <�� S�푸����h �x�������������I��p��z��)K(R�&5�+^+c�XM�����/  ����������u���������	���%s:��	�Ǎ� AH>��1��Fb�����Nt���7u�����v% =<���j���o��b� H<WV�^&��� \���$����H�(���0V&�G*�7��P�F
 &8gu�*�(�'ŉO��a@7�va��� �Ȩ����v�#~V�7�PRR������Iy�SQ�w ���%u�O�����4��Qy�W��D�A"AfX��*�}��"�?E�6;U�;���  �����wJ9���F�$+��,�'�y�DSZd1��""������N􉙭��L�ID����@�D�� �B@�ǸG�6丆|���@3�h�b �����~uD��G �;6�+:B	p��9��H�L�3Ɩq%!|���P����F���>������V��� D�� ���@ �W��D�� V�&W���F�tÍ]Tu���
b�n� 8�qm.�� i���u:1�QB�T �4��9���iT ����V�Ҷ-��Lu"ƀ��&8Gr��7}W�ap�R��Dj ��SA�=�f�D��$�iG@�U�,z�k�֞��v��IyA21�S�U�3�f������w�/$?��􋔰��9u�u���;�tJ���#U�
YP)���(>I�#R������� i�`g6�	O��Pg^����@S`P��?�%�o��6ҍF!C�`
� ��)+�䷉�jClF&A�LL�xt��z��y�����&�U�H�V�;�� �P�X�$��ډ`�������0�
�eȉ R��
w�շH�"�<�6����}�\uO�Ƃ �b/cC�%��	�r<ɐ� tLڷ�&��t�= �u3J�L:�:O�g �t2���V���V�� � ��
)�w� 	����#܌W;
���t����������
Vz~�BMa[C� ݲՍ)-)$bj��z�&a ��R����g�U� �v|-w�w ��� ��I2� �'��$R%� ��?Xx�l=I��|
��tv�=uo��^X��@tt�u"�&������(U�t5�� 5�|��(ߺ�]OF�v�S���&�`�q���4�XR�w��` ��uL(� ��΄�� 
��@ ^)��~3 0����&��o��a����� `�`�o�D����%����{��������{����El�P��:&���Ǽ��z{|��}���~6�
�/�ǈV��
���w��L���>�����U�"$�N"�D���D�^x"�&ri�U��*8�L*t��SW*�*�!�*ȍ�vv����%���Sy &��N&�&���&��&&�N�&�:u&�&���&�&��&�:Q0�L�j%&�&u�(!�xF��;�]
 � *3�!����vj���� � ����p�&�% =U���P�����઩�Ԛ�������������������������T�sM��g�H[�x�+  �= w����.��V��  �������� �(4�Z!�~+���duZ �l��U��]��<���^���&��zp^X=� t5-x~�u:�$f������&����ې- tѐ��t��(��~�u@��z^]�{�9 <i�!|�\6�~��j}�E�n�@fk-����:�7��o� ��'���,�,�ލ,�,��Ҋ���F链�(�i�(�(k(
e��jj�z@5}z�*A7}R�)7��\1��ԍ��� �i�暦���i�����i��������i� ���ڡ���si��e�i�W� 2I�HH= wA :��.	l	�	�	� @	�	
6
^
�
�
� �
�
�
�
�
�
 �(8HVdr�N ��
 }(���  Fn������"�(��!�rg�"�> t
!���'#uY%sI�F���� +xFQ���KQ������9&u��JWǿg57�����Ƈ<`B��o)(�JP��P�'�~_�6���r�^-�؉p^��F�"���F�t�G�jgS9ZTh���z��u	�~�
)Vny�Z%*�V̕����V�wg��v������&�y�ou/by(�UO�#t�o;x$��[T�]=u)wDĎ�Cv�D �Yv@�wS[��V���W(vx.�vK��+N�͐9�S��,�4b܀:uFI�PD���1  ��n-A @@��N�QP��2��;v�t�Uq]AJjV�M(b��tc�.uLɠฤ�)E���y�B�,�z�:��PRZ����Y�k���N
-A��>��,�N,,�,�N,���,3�,�,�f:, ,�,��t,@,b,���,�,6,���,�
t,�,�� ��²,�Sf�,�),�,�,�, u�,�,@,e�$�����o��u��t`-z���t�N,��,,",�i�,,��iF,,�,(��� �,6N3,	,r,�fB,
,F:`,���,,X��,��J,L�,�,T,�N,�,,3:,j,^��TT�h�D,uJ�r,T��z,Du؄JT,؈�D,uJؔ,T'ؠ,Au ئT, ج'A, uJT�,uJ,�,uJ,�,uR,�, ( شH����!�〇 ��� r r�� S[�P��I	� �VW���saCPWU��3��[� ˋF
A���4Z_� S2�G�[3��Ҁ)� �	t�?XR����X_^��>�.��A �.�>P.�R�� �-��r���r��&�v �QW�����_�� �6T6�VZ� #ʃ����XZ��vB� �a�&� ����
� ����2��| �)6�g y��� ��� �r$����C3��� �<u�!r� 
�='���r�t�\�|��<N� ��{""�t�=m0��{
�8�>A��Q]f� �T�U|��N�)� _u���A Ͼ�J� �/f �>� D�LNct���".��� �PkX���0�	.���=:\u-G����� � �{ ��<.t�	��������!`!����øD�<��@L������I�`� ZC �'LMDtA� ~3��Hf �JDF�� 
 ��t���	��� p�2���@���!�R����	��>�� ��裏#"$����BDH���WD����Y D�_���t#7L��$#Z#^�x�� �ø B3�3��q��?�@ �đ
� �� ��H�&ώ�������.0֘���Ɗ1@P���6-D ��X- �� +R����1�HH�AJ-��3�	�(`��&�l� (o��nq2�� 0��.�� ���*��;�r= ������2�����
 t `t�ðÃ>� ��t��>�u�>�I16u�0���u�%�%ѡ����uȡ���	��t�=z��M��SDSP6.0BL G� w>��2 ̏���PQ�Pp� � r#�Ɛ�WQ� ��Y_t�� ����YX@�������&�E�����  ;��2���� ��� á+ �U�F
s?�j�]m�o���=	LN� ��3�����6 wr�Z�Q� � 0���� ��Y���"X��
��>% t���f `d���;�r��� ��R�bd�o�I/<!�[�xIYr;�	i1�p�h@�fE1��lVn93;�f8���sV�v�a߶�Nls[\Q�^�=Y�o�-c�1;�s_��$� ����^�����6	ܮ�=v�L.��jr6y� l ۋӡ6�1;������p����B����P���Y��s�mH3ҹ ���fp�@�3�VQp����2 �%`��ʋ��R 8�P
�� ���u.���+��� ��� �t�QV�  ^Y0v��Y^F✯>�Q�OY ��݋ڱ�����CP.���.Hp.�J���.w�r9d�r\.y<�
RPR �.ZXsB������v .;^s(. �6��PSQR�' Z�HY[X��uB�"r�@Ku�Î�xl~��l�,-�Y3@�ظ���&�tח"D�F&	�h)�;�pth�I���$�����j�1��F���r�P��=i.�S�&k\Cxچ�[��l��n� L������[�oğ�S�v<:9�ԡ,[;vrud�1FNMH��HÌ�	 ���?��V2�X��!V3#�33%�'�33)�+�33-J�BS�3�T�Q��U* �X�,A�[�� �����
�g��,Т \�]�,^� 8�/���$ �{
����T�vt����'��"�� �/bx�
;s��9�|��egN1gB	�[���^��&�GǩW���#��� �H;�|'e`p(�? �r1��m���!\']vC�R/5�+q�S&���x\\ = r���+�� ���Á>����+���9*S�Mr�f,�G��	��d(s7��#����蜁�; �6PP  �C;�uP��@�3 X��$�c���%��.7#�$�3�g3R���h[�;ft;%�* ���ã�ԩ�������� ʹ����%X�<a�9r<zw$�c�g jA�s�I���F�AT160�� ������� 	���fF�������'� �	,�@�2���Ϡ��� ��9Ę�g�J������6�Ȏ�� �.��t'���s���2��Zh�Y� L�Lk�w@xejcc��{��[�oL@�&C"L"��(�<��x-��D����Q�����C�'�aĉ)�cRB,^s���?.@�� ����+�@��U��j�������#u�����ӛp�VW�- 0���^� � �
 �F���  �F��
�N %@ ޛ����-�@�s��/_^]� �v�TW�]��mb0{�b2m( *g�4 &�=DS�u#���G �`[#�.7[4[
[U�[3ɩ�` ı �>P�mt&�_�}^jQP�}��*X�[���R����/5�!l �%�J�RM  �IC�/��CIu��MRu���>�y�[�f�L�B���J&�J�J�^JJsTJ���J&��>�. ������� ��0'+ǉ}'`��&�C))Eff
��U*�߃��� @�>C9t���
 6���u��?��VO` *&�f�.�� � u�R��� �p�r��[9?0q,.�).��.s0lZ.�&6���   ��SQ�CJЁ�P� �;�Xu����+�FPH� HZ�ܲ� �d�>nd%�z6/����?� � t���[�d��u�A �u���u�:<E�[.+=��u��?��P{���((ב� , $�pr�y҄��I��a ���%�%�D �s
F�a� �z N�~ u��q
$������%N �C�
 6?�
hU�W��:.l��L�x� ���V
�^�F�@$� r��5�<�N4q��A	�Q�R}� =u}ib}`2}])O�X�IXLX�OX�9 ��&Z� \��ڎҼ�� �������=@p��=���v3t�������q �0 r6V�4�� �	 �� ��%��%�t��x'� 0^;|s�|�>�%�7�@npWEËD
 z%�б	����|`�&�JME jT��Jr�t�a �VR<0,��d��@��%4��3ɭ=�8u��6x�%r���+un);�t� q��>l �.x �v�  ��t	�s�Ī�6+>h àH�VW��2��'�)# �f �6d �j(qrn �6 N�����tnƋ���6��*�%�p-@��_^q�����~�3a/� �L�&r ��`�.p4�r&�&  ���hu�`� ��ˇې�� ��b;` ;t�h���][v�NڵA4k�'�u��:Gu���uu2�`0�s�m������ �����E�ֈu�������(PF�I�A��w�"��������+�Q?s�S��G����م  m��tNA+�S  ��S���r&�PIu���/� �P� ܍�.r ��Y���1��^ 
�y  Xz����s%ۋ�*� x��ƀ�6&��  �̀���À��"�í'�	yY)$,Xx���@s)V�W��6]p6�a�@ �s.��@2��44<;�4-�.�]//?�g w�h,��| � B�4*����5����?s*C�@�� w=d�d�d��/Hw/@ /=/�x��Q� //���^/A/I+ҋ�h����O�%�L����������$��/�v�;lǆY[��Ah t ;rX� ����QW ~���d�` D��EYE 
PIu��p h  _YÎ�Y�7�(��t� �Ã�6��%C��[.������ғ�u�+� �˽ �  ��!�4��u�  �Mx�������u<�΀u���?��5�u�@2���@�������!���p�K��Ȫ�?�'M�����$��b������^^`CQ@�Td�dd+d�%������ȃ�\��k�kZ��oZQ�XooݾIoko�!ooD� �
oo%U��ooyo&�
Z�Too��oko T�ooɤZo@oM�o�o�o+�oo��'
�]Zo��ooyykA\\	�oO��(Bo�m�% �+mmA�m/�	X.�m m�4miJK�Zm���u��_��	"M_v�yjv���vD	aR�v@vN�vrKc���w^�Zw� ��
wu)O?A�w0��b>w`��<���mH^��
r��C�o�r��o���o�L&o^o�  �����t��?t� �t��xދ΋�+�&� ������+� ��ڨt&����j�+�x���1�����@E���t#D��**�'P**��t1�u'
�s'�'��	�`����a�2���\5D;��88���8�/�J����L�=�x�� ��N���1U;�#�yU ���4�e���	H����� u2���/�����7������^�/���x�u���N#� �^�8��4�Ӝ�\�:��Z��������H /�[��>��i�����1*�*T���kΒ-A����4��������Ȥ:���Z�}�/���������g�,J��i� �}�j�6�&�'�����4���4N�R��S���	�d��9��x�/����� \O����B�r�
�U�T��)�QOh������>�&�D�� ���v4���������,���
i��r���U��@x����y��\��N���U���E�&�����$�.���4�����4��;��S���u���/�� ��� �!! �����|����_��)ڮ��ܧ�V�GU;�&Ӊ����4�`������ x�9t/9���N��7 ��-�Q��ـ��  ����sX% "����I <ZЀ ��rF����� dsN�¯Y�C\
%?\B\0�% � <c
�ܴ  녅�u
6��%t
�R�<�
u��c� ϴ0�!<s3�P  ˿u2�6 +��� r ���ׁ�n��s����'P���Lq7�Ɵ�H6  ������6����6�gxD���P
��o�&����l]��+��۴J@ �2����V��p�+� \�f�"���њ��0&�n3���6���#��݊�>�Ŕ� �.�V I 6����� 2�6�>$`����uX��(��߆2	$� � [x��������%�ۋ� �6�.���&�6, �8���3�a�4�s0� ��6<��rr..�>��3��= t `4� ����t�� ��u!��b��� D���,Ar���`n
ª��I�3s����D�l
�t�� �@Ky�@��� h�	D	� �r3���<� �VW���
Q
�`lu�b���9�6�H9x ���*��Hc 	Z �J7}*X
�P �u�~ u�F��s� u�#~�	_$�^]�/�  p
��� K�>� t������; ��s���Et���
�5�� WV�vV������FP�v
�6�:��F�3_��0��^_���@@Uu�P�y?
4i?k:BE���ED8^;Ǌr$	�3*�D �tH�Ʒ�ѸB��K�u�mFV
y�y*��6�V�\�$_$�N��nV�K�3&�

�=�
�F��� z�׋��~3���`R��u�
 3��+����؎Q�K�F����I_���P��]�F�v
�����0�LAs�X��V��6rw�3t����,) 6G*�$I���WV��O��M��9b��A+l�ٕI|�����z^_<�/��
�tpJ���2���)�GD*"'��mA��MV�~ X=��D�3�&:�QE�wtII����; �+  ��V�㊋动ܮ�tn2�Ftf")�<$� `��^�&�G&tJ&�
T	�7;�~@1�&�8=u%V�<S��!
��u`@W�@�
���r�+��^��ڍ�
��t� 	S��&�[��!�R ����(��u��]�.�-��WV�6�BG #g�2��4���A,�TA0����Q�����x��.�&� �؈�V�$tǆ$@DujiBio�>i@i8~�i<ia��j<jM'/j8jV W���]�M�Uu�u
���]_�!�f�E
��)�f)�)�)
r3�`�E � L_d���D"�Yy  �+Џҏ�#��z	f ��� ��u��A����>ԏ t3��#&#�#1#�a�4�<  �=�؉^��F�&�G�
�J�J��V�*O� ��,ϊ�P�C��PP;�Xt�<u�Ӌ��� ��Q� $ �U�~Fne��W�j%^�Nf
�쎋�3܎
����"�?&���-%�91<���F�N�Q� u������M+M��?�(��Q�Q�@"�DpS=z1}w�,<��,�<< ��� ,$)<&,Y�y}�\~�#�n8�t?t�\s��n�N�Լ@\@����;.��� ���F��V��RP�����#��
 &�o9�" ��5�88bú�+���/v6�vcn�\N( \Q��? C{[ 
|���  D���V�w�##	��� 5�������݉N�D��q�� @P���� ����C���!	��5J�
������w7�@�&ݤw�s�T@E�(���$H��&9|s�D��j��Gq�)ج<���;V�e��N�-��*��D������|
�%4d�R����SP���	 ��N�w�S����g�CI��C����2؏֏�� �%��+��z�$�v&�< t$]�"��8�7&��F
&�AP�? u�72!�^V���!&9v@M
�
"��0M��_��Y��N�v��MR�$e)�&��rPcVwDvz��t�d�
�nS�x!��&��a䭋���:?/�/QPS+t��K-4JJ,�z/ﱓ���w� =�DcOp��-��n/�U�o��~��+\R�Ja4|�?���P�"�A�يF\
���&8t *3��ǋǌ�_NH ��G.0�� x-�&�'C:�t�,A< �ɀ� �A��
�:�t����Z�����rOs�
GQr���t�%bȌ���p���,aVsQ��C�u"��$�� �0���ЎYB G�~�����Ȱ�ҷ��C�� �3Ҭ%� zt"tX��D�[�
�/�	�IOWV ���H����+�۠	#��@�+  ��u���u��  ���uˌ���IF�&^_�=RZX��HW��JZ��^��^�^���g_H0^�8�V�`�t+�L�ч��
���Q�7�Q���Á�U�D�_�K`X$u��x{	d�B�P���|�^ p&� t���P�(�/K=-d� ���E�4�9j��i� r�����sr-.K͌pj?ig�dlU":� �G������/t\t�:t�\�.~G�#���	���כ�t��t�t���p�
�q��V*C5 �r�F
t	���w ���ܴ9��';+(��t�d�: ps�= u꒓�C�R
<?=<*u�k����@�#�/�z��.����҆�C�V���o�v%$�J@R���	�=�:
\
�<�F�G&�F���W2���X��p! � E��Q��2�5����"��أŊ�x�t����������� "�V�u/9`v�~��V�  �%P��P�*�"
/"� �^*P��^+X'G��V� [_�p��$Akab.^^H�`.�r��P78��O>R�A�[C��<A�t�Ds
=P �C�ua��_��<#�	�
�d��O9�	��N�/nB�.NuiS�P�P5�D�ڋ�X�X��n|JiQ�
���2��=Ƀ��?�OZ@���&(OVE�00`��T�Q3��$"�{�7:�A6=$ ��u� �g VZ�D�\�r�L�^DB�
IF^��� �+��O�w�ʈ�G*��@� x1�,aF0�/�O/w5W��0S����+7�� 9�߳[]�|�" ۹�"��)��.sA�VS3���X}G�������yR�
�ԡ�?O73���؆�d��8�������������u���f���``��r;#wr;l'vND�Ou_p}c�� [�ĺEN<Q��Ru	b�|SpR(O��[	H2S�40�y������ V�O�j^��ѩ�ۼɼ�)��^{O�_�N]��E_q��_
"�]]+rVLe��S��5~��=�|����6>~nmd�9 �B��0&�������HSQV�*K�H;�~�I���_$�^Y[2,0'�򎿔WY�c�$�H���:S��>ߐ��
���4�7 z��V3��B 2���2�q�����Ut!����4)~�L���f��<�ut)' �, ��3��� �3�9�u�GG�>�b�^�ѿ�60�� �' p�< t�<	t�<to	�kGN�{�\X<" �t$<\tB��3�A<p���Ӌ�hѨu���91+1'�\O1�1u0�1����݊�G��B��  �+�ģߊ�ኋ�� `6�?6�W���6\"�����6>ӹ���*��u9�f!�~�8���"ҟb���^�'���0��\����ժsL�"��.�\4*!�4��J4�4�/�4͔�:�G�.
���6��, �ÌF��(3�3����t�>>oP�F�� �@$�F�����	 � �RP�����㊉f�dV��ϋ� B_I�3�6;��uG���p ��t�^0��?�G��B���T}N�W@׾���;�t@�t�Q@x���떒I����f��"��X� ���nk��sn^�@ˑ�6 r9�Ks�P� X2�L� �=��� ˢŊf �"�>r <"s r��<v ����ט���Ê�����W�v� �D
��tj�@uf�Dn[ݑ�9'Y��� $�$�#�������|3ۊ\!uQ��;u�uHmf����$�u&���t�Q���~WS���	Fn��L
 �eS�"Tn�[��atыAT+�B ���UJ�T�%QQ�tk/�Ad��AY�|,M�;�u�3�K,\�"ip t�?�P,��,@15���_EHx��&�!���*��	�.�T�X�-ʍ��C`���t!�D��M0�'Emp
��V�S�$�P| q[[�t�J�Ȇ�Á��ft- L-!�
V��y�a�~_�8��O$dqD|D H �����Dvqخ:�`3 �o�F��v
&����~P�.  }g���  2�, <Xw�$�� �x��2�����:p7������*8��V���6�(�W��ȧF�k  �0e�뛊]�6<-u�N@���<+
�< uR
�y�<#x ��n��g��N�� ��*u�\�y��n>"02�<��
 ���k��F;�k��UD34�(4Ǻ=1�:D1��
��)Hl��"<F�
 ��
�<L
��q���N!2d��<i�y�<u��X�x��o�c8t<s�ntQ< Wpt`<Et<G ���� �������O7����p/�����������uW�N��2�rOY+�����8p.b���뀢R3���;��0u�2�9�6 ��u0�F�ufR3�o����y���XE��Ɔ��:����Qj0/�/���/��M�F���$@ Ѐ�~� t��P��P
=g&�Y�/�v� k�VW ��t
����F
&��
�
��!���tMu	/����gu_�������-�eG���W� �� �����]5��K'\��� �0�QV��V�i'������L���� @t�� 3��}^�w�� ��Hz�}�Df�������p� �~몊N�sv��@�t���0tO&�0A�ܟb1�?�-;L�� +�s���K� ��+�+
}���WQ��Ȳ �l � Pw|�N�� ��Xt� 0� Y_P�v�t5� � �`R�v&���	&>���' p;t������������`���Ø}�-3�Oxn�?�&�G����QRSK\>��O��ZY ��������N�W Q���������_t3�!��z���\�W��
q�8�l��Ɠ p���0<9vF�7��N��Y+�G���$ W��!P���3۸�P<-�+u�9w,0r
b`ҋˋ��������X-���;;� �Y��� ���wr��? �s�~���@�3��RPvr(김`l����SQ3�	R?���~��n��'D
@pN��+����	p+��L�v�V���͕�~� }*�P�v�Re@�[�"f&Q�v��g`�L
�ѐ� ����$"���H~�;��N��� �h��^��l
l�Qe��R������Q5��0��@5�D�����\���~�\&9|�u�+z����T�< �+$G�SQ�z�Y��\*)~:)i�a�b#�<m�ܮ_F�-�c��+.�T��  �ƌ�N��>D���^�V7�U~:��V�ď돉�� 0ި���� q3�D���6�6֏����3�U�%���2�G��Џ�nܔ+���XM8�\�&��� pJ��ٌu���'F��|�G�#m�o�W�o�o���)����@�ԏ6&�o Pj��}�� 
	~I�
�
~
���w
�ƀ�l���~um�_����h��U
j�8���$<��w=��F�ƹ���эD�����+ �Ȕh+V� @�e&;W|	u �|�< ���|�u4|�+�^:n&WV#l�D�n�nt��V��W��f�����s~G�'F��o�BS�p���3�1��i"�D	y�W;=@Aڙ�ӫ>��u0����K��P�_~����Kd/��h{�F��^�	�n��X^���:�;Xld�V����t=p�Q�#}+;t%y%�]q�v#u�4�.�-��4.�+��$!90N!u9#u_��s� �+� @��a�J��%>:Fg\�u@:2��0PG���ɾ{o�VF��t�G V9��=��e��T%u����W��. ��?}��������(�	.t�6�'tV<^��	etE�$�$�ÌT���N��0t�ǝR���^���� '�<��8���9����f��r�k�)�q��EHtA dGK���-��fE������ r8bMV��?X
;�>�����~��F,�
q�> � t9�F��]���Q vp���V���V� ��~ ~r����<"�[����&T��73��F���;V�13��iN��qm��'F3ˋ�`}Q�h0
�m-Rs��U���AyC;OA<��P�ef���W�G���Z�T?�8?4E�ɒd��\�S��8ANy�؋���'-'��d|i4"( �T��
��
�icڢ��ʸ���vA@TM�W� W@*�@�� CH5 �"�9Nu]5��� B0�C��J	�p��G9P��اr7H��A �̗J������"0��!�ih��aU�&�&���G}@ �	5������	;�X���9�B?�@%T�0 ���h��4=��}�}퐺6��H���H�"���~> C�b�B5K�;9~ ��*��$�����J=��|�|�$��32���>1 t�T����;0�G� 5"�T~e�x�Eu^i;a)����)�;#fu g�;��ސ9���bO�%���@x�����FHnZ46  � ZZ�u2��*�P-� ��D��"	 ��&��>��O.a�$ݸ� �(9�	�e���2����� �= }d�ɍF�P�	�\����z����
���N���uӍV�{����_
���y����$�)�GZ"2�I.�@��;�)���SK�Nʠu� u��THTy��]�E"eH\��ċ=��׵	-v*+=�|����0�x�>t�g	�S�f�SW��&1	h�!e�rµS�P	���Z�D�R ���N�O ��F����CO(�~R�;�T`��3�(�����õ��"�Btk Z0�-H릠�p�+a���/�
,{���|�&wv��w@���]�l���c /w*�b/�g3��~��L�91}=�aHP(����}W+6:�f��3�M��E)F������*Q�"��.YZ��+س J�r��RQ��F� @u3����.SQ�b� �Qe ��Y���t�d[Ë��л�
	�� ށ�����V��
�{�� �ڍnG����=�&�Y�F�"WV+@H�Fup�Xp �_�v W��$<u?\����2�h��ht-�+V@�F��~!P��L*�H�Q��1�9;t&����]+�Ez ��N�e�U��\�`��~��o ��8��96Ԍnrуt�H2V��0R@p�t�G���u9�M��ZFR��LW�);Ǌ2�� 	���vd�; l�B3ɋ��D !r��t|�^��F��
�͉1���+����f��pd�?�
��Q�'���w=� vJ���ܺ =(s�� ]���5 2�<
t;�t����`�& �y�u� �N`K���� �R�m����X8��PSb���+��Q�HYr�;�w0Y[X^ßw�� �~� u%�s�	�$Cl7�
�
�?j��9��� ����/+�E�l��p$4�uSw����fR'^L�r(��M��&� J�J� �7��C�ђp�(u�APjE@�j��Bl �J��������Z�ڲ��SxF�$W�~(B�Fd�s�&���@L�yεO��L/\P���N
�~
 �h$o|285|������@�D9t�&�q�1u
��G)4ކ�K@�SJ龦S��
&� 3�����[����	
iT�b��&��Y��^�V���F��#NWV�ưV�v �D~VW��9��T�xW+� �sPI�s���E ���� @�A��H+��#��+Ɗ�@�4�����E�\���u6-6�[�8�7����8����+)��4��@�lP��ED�u�Cy7�I�y� �c^_]ˊ*�C��/O(��S���? �<w�7� �
��[n_�
7��}G ����� $�����n
�
��X$���OyC�W�H�V9D����í%��"��f�
g�r;!w��%v+F
V��Ch
��� _[��̜j�?
�����_3�����e~ "6�E �Āt���f-%����ƴˋ�aFtM�e=Q�u`0�u���= ;`0
���6�}�;?t���� �$����5�}3ɊA�dy{�  }�m
 �\� �~���M�� x�M���װ��� 0������CW�ߍ�$PW�,_��~�?rG�76�������u�F*t�y ;�= v�\��ܸ-�?���1^�D�v
�n	� 0����������u�ͷn��� ��	2��^�N�V �v
�f	����ѷ�1�������%+17��= "0�KW�l -u�ilv��<5��r*�L�'�9u*O;�v�G
6�&� +���C6�\�����	�0�����&�AL��A �����؎��܍v���6�� �U��]����Ȭ��	 R����2����U�M�E�]�ڲ#��M ��F�P��,N�Qh|�����7n�$ bYZ�J���;����E�u3���QW�E tf�� ����/+�IA A�w�tO�s	'��5���3�B�
8�&��r t� ��;�rOu�  �"��r���H���ws���#�R`�. Zs�t���� +W��VG� J�B����_��Y��tJ  �N;�r9W�s6BSQ�� ��Ʊ��u�  $
Ƌ��+Î6ش�J[r��6X8����WI;[70�=gtv�$������OO��_��+F�t��F֓Q� �Hi�f���?�߾А�0����@� í�/��t�$��t��.���������0�����ĐWV ��^�L�dfE�D Rt��y�-���l ��S�5>���f=P����X.�9��7<3�@��ː����
 ��~�
��9_�<0�/�4�H>�\� )��AtG��9:�"�W\jy� ;���������J�8�ً��� ����������֚ ���ٿѐ8�2�QSRUVP�If���f&u�`fY�Y���iُ20��OI��K��s�PIZ[� E��@�&u��Q@�P�G$������ �����4��  ����N@ �p+���  �i@�]�%��O�@q  �וC�)��@���D� ������@�<զ��Ix =@o�����G���A  ��kU'9��p�|B�ݎ�  ����~�QC��v���)/  ��&D(�������D  ������Jz��Ee�Ǒ  ����Feu��u  v�HMXB䧓9;5���S  M��]=�];���Z�]��  � �T��7a���Z��%]  ���g����'���]݀n �Lɛ� �R`�%u��A �q=
ףp �?Zd;�O��n��  ?��,e�X���?�#  �GG�ŧ�?@��il�  �7��?3=�Bz�Ք���  ?����a�w̫�?/L[  �Mľ����?��S;uD�  ���?�g��9E��ϔ  ?$#�⼺;1a�z?aUY  �~�S|�_?��/��� ��D$?��9�'��  *?}���d|F��U>c{  �#Tw����=��:zc  %C1��<!��8�G�� �  �;܈X��ㆦ;Ƅ  EB��u7�.:3q�#�  2�I�Z9����Wڥ���  �2�h��R�DY�,%I  �-64OS��k%�Y���  �}�����ZW�<�P� `"NKeb�����} $.ޟ���ݦ�
 �VW�~�
;�  tzy�f<���F��>L�uaQ��>�5���=8s+�n�`lW_��T;#��"���W% t�S��y ��2���fH��[��R�7��pA�A|&�m�]_���<�o����.�w
�.�Osh�ѐu�QP��\��P� U��l�T5p�չ	 ����~�3���)ċ��Dv�]D3 ˁ�H�N���#�;st�#�;�t�7��Ӂ���w��?v�"�B;	.1t��BH��&E ����?�T
�ǀ=� �^�Q�(� $66W6�W������YD0����u֋����V��N�^q�W��|�*�_�f�"�����ئtM�y�׀��rw������[�  ��� s����D�sV�|8c�\�L�X�	@pR����wݳ�Fu��;t��N����}RsFDFD=.�뾸_���U�]
4F�d�v 3��^��v�	��@�m�F�� ~̬< t��<	t���<�t�,���<+t	<(� *��%0r<9v<.u��w�~��=1N��]�5��N�g���f=���+0!0[,0��u�")�Q�-.t�&z!;**��*�-�
{��^惶�\  ��^�3�<Et<et
<D Mt<dt�R��D���8?L;-0Do ��$  �Z��fw����:�y��?f3�^�+^�Ҧ�P�H� �Ov&�p��O<r������z�O���F�����P�{��/*=P|U�0~ =��� &&�v����>ܩ��N��"��(���re�`es�̀��i��v���dU5 m
������tA�v�r�Dn\)�u�o�*�"�VN�	��~3�9�<ޫ����'�Kj��@�T�o�2i���¸Z�)����02���f�T��R���H=t�t��.S���Ц[h҄Z�h���F�ʅFȨ���J�F�h���Fh��F�h���Fh��F�h��4Fh2�F0h�.,Fh*�F(h�&$Fh"�F h�Fh�Fh�Fh���B����C��W_��F �.a'N�a�S/_a2T![��ú����D�vf�;��pYȋ�&�F�:s���F�^��Nˀ���{ �x 	��!�f &��-�� BX���N@��RËً�3҃���x���¦N��
�6�D
6�\~D\�@�L�ƌ�Ś���6�����P5���$����D^����\H�^�K
<��E�Z�w�
@��� ��t� 	iu�'\9�m�/ �MSEM87 gfw.  GW\ ����  )n�V����w��.�7.��p+  �T����NOC=
�V.w|!͋�

� 
�r��3u���e �U �t��2���t��P� �O��&�
�t8���O+��ϋ������SWQ	wW@"
n�Z WT��S[�E`Y���>Â�B��Q�	��Y�JR�X �>��&?�?uM�@����tH�L��hjj ��'��>_t  ]
�*%s�����j0�h�+"'9&� �@�13uj"�"9�"�D �2�]�fv��Hø�6t����ܧ �6��H�Hy���$����6VF7F�s�E��: ��C��� ��]�^ùb45�  ~�!@��E������E�(H	� 3���+/%��/�������=H%H^��@G��3�\�A(�bܛ6�7/6�G<��F������ ���tB�+ )�������9��� K� ����C�PU[���v�����F �FS 7��(sކ�S�~�&%���S�3��,2��>a�����u
n� ��m��u��t�����''���9���������"��z?P�0p��=�OX��3 %8= Xu� 4��n 	  [��]���X�PS���6�G[X���VSQRW	 ��N�ӊ̀�8�p���˄�tR�����u�a �� n@u0��4���t`t	�'�   ���?�6 ;6���~���1���<�K��4��J�Z=:5����� �B�+�D�f���@��L@,�^Z�:�ZQuP������%>J �8���y���.O��@�-<t#��OR���U	�JU�����FF������P��y� {����ʋ�����$u$�0��_���z�À��F �f _ZY[^�gF�� ��� Q�NY�� ���tm��8����t�0�0uT��aG��wa;Qj������� �^ Y�NYM=�HM.��^��9� �;m؛��(n

 ���:$���@Mɛ����>c�n
Y$��-�0 ~�F���t!� )F�u��n���~��>@6�"�3�z3�C ���% ���=� Xs| �������@u\Γ�QS���)x��>V � p�ـ���؀����<�E���`��~�~c3_��F�c����^[YM0���S��f0`u8��u1���0�+��u$��� ��� ���u�� 0�u��� u����� �� s��L�!�@[�Xϣ %<��8Q�3�.�
v����-���$?D1��(9% � 5>2�������G�L= Q
�& U���]��g�OE)E�:C
��� Nd]�Ӵ� #���#i�#3�	��) �ъ.��C��C?
�  �tّ����PU�V�������Nq�� ��$&�İ��.�S\�  R-�=��2\M83)#3�  TX;�u(�@%�0=�0u��@<�r��=���=  ��t��[^]Xϐ\ <@�ZBRx�2P0��dH�F�`�"�?�D����$.&	0:= [eo���  {������  0d�h�J( m���� � �  � � � � C%k%X�$�$
�!"&�"O� R b T h o ?��T[v���Y��f]k{)�Y�xt��'� �%� ��_�d T0@B���%��@ ��
@��?��	9���r�" H���j���0�����Se�B׳� #,�k��
�<�@Kd��3��W�E5�h!��"@����Kx�����\);�� )������ �`�y ���r�T��{�Z�>\i��7M�,�x ���2��f�pˑX^���� �2� y��	cfψp�9����F����	�2 2[�ɤP���r����K��� w��+�RJ�� eBPU��� q�K�$��C� p�8V
Ob� m�m�QP�;$��m[ �P�2DZ���t��P��T=�� ���_��J��� &ow{8���
]��{����~�	�H�-�~w���W q�:�O1�5^<����K�z��Ӳ8&�(	/�Ċ}�vX�vp>[�� �R`�3���&���l��_� P8q�v|� ��������϶�!�P�RQS��
 ���Ӌ��~GG�`�M�����  ���.��=�F�
��``������F�W`�0����%2��' �S��Q^ 8P�����(sώ;���$��yF��4��1<��V��T� ���t���p�v ��ӊ�G|b��R���3�b�B��.5|T�.��%�.�n �4pp�5GGN������� ��  �������t
�tP���S��k���S�[� L�����>� ��
P3�.�>I�ߎ�F�V�UK��^zS	C ��� ��L r@�6>��q�G��S��t(�%��	�L�W�����9!��Zr �?��Հ���� ��2�+�;><�����#�]q�[YZ��Z!*�Xϡ)�㜟Њ>���KA
������u��&��p��u�t�2��р�w��qQ�V��J�V���9(�t�t���� �r�H�%G��$ԊmSY�U���*
�
�5P�:v �:��U���
+�
	�B�>��t$��
 u���t����M�k��F�  t�F<	<�	��O��`	S� 0&x�P�u��u��t�s��@Ð�J�#�  ��3һ�	���&���
h�h`E {
D����2u �
2T
�M�D@�'�����Q �U
��2[��?=��	2��� ��R���IX�
�	i(��.�� D�_�;�t��8�  "�2�x�놋Ƌ߃Ƹ�����8��r�����`�~�+�|͆���� �=C ~/UR�u� ��=y�݋ª] 2}S�x�`����� ��� �/Q�*��譋���ح3���
�p��|5tƃʽ�ы�3�M�w�tSr)�|3��� ��Ċ� �֊�͊�ߊ�2T�+wt(��v �Fu��������? �� �5�������΋���� �?�Xx" PL\|s���D��s  3@���+""op"����ӯ������x��'�X��  �P�U��2�R�@P"�n�3ۋ�� ?��t���H��U3��U�^	��ڃ�s�1,&PX�P3�U�2���d2��Ik>II��I�I
�e�\�ʤ�VCZ{V��KV0#Ձ��?\�\�RO�M^=�Ӹz��Q�U�D��}���C �n]���I5}�  �^����2�UR��VW�_^�	��@������ @3��r��q��EU�>` �J W;��@
�<8 �����t�r"�>;Tu;�u; �\u;s���
���Y[v�Q�6� f;�s�b�u;�wA��RS��=��F�@���P����F��衜0�� ��[+� ��[�]蕒��sO1�?7.�{es��O+�� 6 �@��ɐ��N8u a��
+�����4Չ��a(�'X]����� 9&\���� �Ǌ��݊�Ί򗕊��2��"�uxN&"x�t���e��
�
�tD� ����r�&��wr': �t"�XP��r��,���v0�F՜ȵ���Kl��l�� 8sv��;+fXǃL��fr��ٝfD@nz���U� 0ᗉ�M�]�E� �䀈e
�� @}�A�~T�u�E_�� �����X�����z��
p�
満��������%� �w'r6��p�t1�\�g�K�i�Gʷ����'���2��S�(�R�3r"�җ�J
&t�Āu���t���&��������$�ȆĖ�o��bo�ʀ2 ��<�t!< t3�d
,�] 0�t�T��|��4�� @����q�F؀�|���E���� I@H����
�y�뗸�5u�Q�� Ru�\�D�?����� � �R��+� 1D
�L
��u�
$ =� }�=��~�.�0���<�ҋT
R	T
t78��<�<�r,2������t�Ѓ� �2�y	 �������t���ë��,�
�x������}M(��M1.��@r>
�.� 
�8��x)����  멀����M0��0R��=�7���$��
ƋT�����D8��s	����|"L8��ފ�%� �HP�����+8>�r�> ��y��������*=�>��  ��\�L�T�l�\ʊ�i�t
2L���4z"pw=�t=#d�-���$��@����u����M���g�2�,��L��~ۘ�y�,{��hr�)	���f+=96AD�L$����W�  ��«�|
�瀸�
�
��B� �\��� fd������(\Y� Yl��}��~ۊpL����RNxÉ:0t9Pt4�������Ѽ y&EY|��&S��s��'F{r
r�4' ы����d
	 5�
�Ã����z(��
2��
���8�
�*
��AB	t����v	��^�̓�q��tI�IT��G�l���/�ݐ���	z��W���1�A�9Ӹ R(X��X2 �ɈL�π��#߈l
�Y��(X(%�`8f�D�e�R��V�0�Du8u.�L`���*��|�����*� �$
�y��t3�x	_�S�Q�VB>QȠ�pi��t=����������������� f���8����-�,�V� m�.8�A���2�3Ȯ|�u!gf�`�]����`� 3�x���������������M��#�t?���?�	:9���u?lu�����R- ��r��H  ��_�Š)��O���5�?A�|º ��b^3��x��N��H�3���� ����u���s�����?�A��_:��9Zvj}� jP������%l-"��2Ʃ��3�� �����r\���݄SB�����L�W�W6����?��I|a�p6�@}[ �~��t�k�׻��ܟ�0.UBs����.��Ԓ&�5a=D u)u1
�"���E�s`p ����ð2�P�X��)��D
�H�u������i��
 E�ć����rڎ؟�&���U숝w�2�=$��%-�m�?��|"u� �Ol,u�l՛���$��ʙ3�l#'#��ܢ�|��e`
櫧�5���`��l��w�$�$!�Hu��v�!l!J`���~K�|]
�u��.5�48CD4�d
�'	5w�#������R�6��E �$*ȋE��M

ɔ��wp=��=p�?�y	8�>S��\��!�3���8�t\��e
3�0��\��
] 1@	2�xF
���y-�W�;u|�����W	w'e�@_9NDa2A�+փ��$�x�C����x����p�et���MhU�!���A��A�� ����	.ע_��bOFî �`	�l
��x��0�������$
R���ᩋ��y q���sZ�n��%.1��̗��#���t����.�칺�����FF⥴���Fv&v9�@���1�I�t�J-��(���論
���0U��k�3���? ۤ�E+D��� �En }��B�;  Dr%w;\rw;L 0rw;r� �>3c� ��e���� �	�s���Qt�}
 CP�Ń��.t�&�� ������롨�W�MtA!�@w4� ���3���UE�,�8(@'O��'��r�{��,z����ш��r�� ����E��,��s �\��r���	1�K�r����`�ӁSG-�D pD
��u�V�J �E��c�H��ظ��T�@�a� I��E���r��9  R�u����W�s��� ��3������E��
�M@�ȃ�ށݘ�]�MmA�Z��_ ���쾃����C��W�� ��_�:��V�Ɏ�I9&�U ��:�uEVW 	���ʀ�� ��:�u(
�w��g����?/�P;�uƧf�u�aS��Zÿ~�����WVS�r	��H���^.��_�o�vQV���V�V���Y����^5��i.[W���>�-��EYQ3h3>�;;9�;�_�"� VT�& ޜ �^��û�
�]��*�D'�
��"	T$%��%x@� �08��s76(��c��<���` �$���	���W��cu>P �7�����X�Q	�H(Zȏ5�����|$��W��T '��ؿ���E��޶#�V�Zؘ7덑�f
af
]�D �Tp$u��w#CS�z���cNm�E[_S�i [h �t9��y���۹PI���s�W��J�$�!��'!c�f�:��&�T��}���WJy�V�`Ɂ�R���^�������T���^���� � `5�!�r&�t&��&F�%�#v�<x�#xl�PR.�.l�ZXq���v#. �.�>p&Q� ��Y�.��t�����I<  gx:;������,��A��V���k������;��RG����(����������;�(���=��cR��g�;�|������c����;�Ў���������x�:�$�9���N^���	              ( 8 H X h x  ` 0 P p � � � �  0Pp����:��������������;��}�Mm .��1�P�`<�� Xt.�.
��1��0�� ttt�/t*  P�0c�XP�=�1�=.t�=t�@Wt���%�(t'''��''	'A�� 2�'���;�U��.��> 7Q�0������5�!���g�/�1�3�	��ģ /%� 6�4*	<�]˒>bu3b?%�.�9.�
6EQT DAUVW��   ��ܹ͋ 3�6�00��%Y3�6�?u 6�l �6�&�=Z�u.�>=0n�|&�E��GR0_^��^Y<�S.�� u
� t/=
t"�D.�6&�`�E>�[SC�r ��]>���u�'����[L��zN[�Ä�]��� � �D� D�Us�>xt�>t�V �	 ���
������=c�Q�xx�����;���������������;����������w�����������w�������������w�����������w��|����������w���O��"���7�u�L��a��������w�����������w�������������w���� ��MS Run-  Time Library - C  opyright (c) 199 l0, Microsof�rp %s��! D��J%c: +�U u���
�  	  �f�5�鉀�\��
�@DBLSPACE.�lRVE�� 	=/Z-`@/0��V4��"ց~ ERASE��1/��u��j �]�*w=�*� [�x X�u2�lR��g����(�������% & ' �af-( ) �b:H n�T$ F�td�b�
 ��
x   �U �   �D�  ~<�S   BN�u(  �"��(, - . 6���F��" # $f�(�����! �+R�dPC  +�(�	��S,�6.6s��Y�s&�%03u�LSG@�BOLD g`-80.�03d�*
1*L�(;P�5*.70 z�

C=�	6ӳ�RE T��use,"f�Z0F�4�9�@^'�C�6
�<#���   ��FAT1��2 	6 �	COMPRESSED H�/�Q�$ � . "� ..:�  .�DIR)�0FILeCHK�=*B�%04d �l25d�  @��  <	>�	dL�u� 0�ScanDiskMpthedirecto><rivf^dil, at��of
o5�clusters";. vo?�O���3a&	no� Bcompessed��]3$t8�z	invali�.you�T�8T�{).nd�l�os�wJlh&fHmui��fob_m��goi-�\]5c",�O� :b��vUa�۝h��(ar"Z��Wm#!�*hooU�axpaiIr;To�a�T0LfR��e@MD�̏s+c�ntр4ns~i�MXk��z�xm�e�٤u�yUw�h�	>y�1%*�moqC}��f.wo��/ngB�D�5�e���u�N���d �r� N `�ߨalrorTMį}s*f��>namZ+axxR�KwEq��yD�أSCANDISKT�d��� %2�
8� I.0� A2`��LĦsl=kDaff��|
6mpt�s�.�ccD�ful�A,Y�17som��DOSi0gun�a�9�M*h6lgd#EAlMgh`$�Jge���dr;@[g� typ	$x_}Ŕ,��7]W>�Howev��'E�Qd�s���itL�7clWm�1�c1]-�H_eaR�h�H�ctuLFO�+��
bY�2fbODQ��S�o��� [lKdy)i	�us�![�$s��w.

�ryǤ�i!7gna�I T�s	jS9u�<�s��d4�6pue]�A� IFfnishE&6s|�mov*ƀ�� D��t�`=��� ����8dGtj}mb@��C��LritCF�i}sV�*:	I� /QzFh�Am�	���phyY�c&��j;��T�ng�ӝuu	tP�sȉuumuGy\DpyǠ&�en�� ��_�
�V��SURF��2S�H�ܮ��#J�St�� ��
gra�i*.|n��J$#m�a��B�<QWV�ny��8itsT�kd鱪�4��?�H��ab��rT��i��rA0s@xlh�֊[wor	%kd�@�s�?}�Iz��{���jr6r\����
uZÆ��LS�m��g<n�N��y-0�m_c�'��z��!s�!s�d@��ify�dR�. ���flop��$�ckupW�_�|kx�ELme�^ Lm%�P0.� 3�p&A&l6r�#�]�CUϤmQ+�B�an�X3un��k��$%oT��M���G-gn����o�%:�d"nnEyt��ص��Q.D�����HECKONLY"ir=�(�7Sqt�sub	�UMDBPB� R�/�8wzNDm�l�ex|p�9t����t&��QX#�&�Z��axis!%
�1}-H�tcr%�de[��B*�BF���i� quiWP�w��uC3�B WUb"B�z���"3�G�Wƅ� 7dx���m���fEJ�� Vt��gniz4��g�m��"�'�e$ lappea;Q̒agm�����Y-DeK
`-�tK5A�;��  �$d(`YAUTOFIX2��i�EN��T�?f/dȡ�%Jh���safls!d D,�2�����C�iialo8!a�cifp��>iUm�d�/4J�rDhG�o%2rk���w�$RI �$\�p��4n  �"�/�Qt�-��Iy�i[Ⴁ<oc:\%b2�e�D�x
@�D�c��l��k֏�"�{��Bad\����%7�p�%���dYH�r�H�rdd�t�RE@@ADME ).�c�b�5�?�w@� '�IH�=<'�.py\xA3)E?,a��#�!n�	�AaH$) QKX� %)=�)�&4.�4�%�w<v$�]�~�ۂ�i�+\I���5 dud�eIM�]��a�dB:�����^_P�2wF��w�B8ύϼ"��:�ex	pTN*�>2X�isrrAm�&H�s�H��5���N%�a"��iZ0\hQ/��S�䰴��$�fuN�af_B-G��(RATIO	S�6NExN�$�3�� ha�;N�LLL�tr�laSB
r�m9�fTYrDD�TXT&�yB�xXԕ�L��$M��C[����iNOSAVE$'��P� OP��ocia1�r����>cISp�a'd>�U=� �,�i~u6֒52�s{rtV�SxB��ac�8&��Eg�1�"5Rh�un���d�e5sul@*���A�S������Y,�_t��UNDO�$��]`Į�K-<��I��mEt�LDܻr1��5�D��� P��eme�?�V��C��P�AeT�Em�dYSIʛƃd,�!ˣZ�"���5Bde�t�beI� j�xLp�-�K45{+�H�hlDNmd�]l)�$o�}��2�rdwB%pRepe_(qr���cm/C2SdXwd8��eemLI>R�߮�wn Z^�b��n�c�� ��vOn0Y�.�W>tO��ys2���$M�olw��G~�3Ml��!!�I��X+ԙ�]t�	�%4`)��x��vP��ndsY�i�ڠ�Y	�20Qet���.r�	0li$'�}T�3	����3b�ltJ��ye� 4�&d,'��P�f��Sv9�	�,�]݁9a
�xPʔsu!0\�" CVFv�$\��t�B@��<�`C@�O6*rƼG�H*�s]Rׅ�o��Uxpf�dwE�� ���+@&�d�of�$-�ƺ�\BK��L�� D
��iВ*�E:FeEx�pt��:,�le>�20,\�7 ��y hidd�&ASSIGW LDEFRAG٠��BTf�t`.ks|�s~�h/�-Ls$Log%��OUNTkn$(�sD����M�4h\�a$I���h��Ҡ�sc��� �:DS �q2
6.���o�
e�"aXw�--&��ol`���Sj��P
USTdwOM b<q@z%H�(SU�B�aH��Ap"=HPFS�UQB6
:e# me*{��	.$so�l��C� = �hel��p0�d��]���U�vi�O�I;hf��m�)ENTER�Bp�A�l~�)��X�AO!�LSkip2�/ J�W�"l�k�eI�p���30TY7HPoV%�x.T$I9T'��.�$�'X'��oa�=(�N�S�u0Ycϴ�ĉ uf#'	:v/�w���p�p@NOG�� [/������H��FS�$s Y��j. (NH�32�[�'���\��n |��&Jh��lxB�� u�qgI	sPCv����
u2${�+14��:>B�{HRX�\dhn��w|�{����������{�������������{������{"'�,1:?��ELT{�Zbf��py�{���､��������{���������y�
�!'-��25;{�BJR��[ek�{uz�ｇ��������{���ǽ�����{���ϼ�
	��"){�.3@��FNV�{`in�sy������{����������{���ϼ�
��{�'1:��AHQ�{T\g�kry������{����������{������������{� ��'-1�{9AJ�S[dm��sy�{����������{�������������{���(&+��.5>{�HRX��^ht�{���ｙ��������{���ӽ�����{������$-��8A�{LWe�lq{������{����������{�����������{��$)2;��DMV{�_ep��w���{���ｬ��������{��� ὀ��#+{�3;C��MWa�{kuyｃ��������{���ݽ�����y��&/��8AN{�W^e��rw~�{���｟��������{����=��`��"{�*2:��BFN�{V^i�t�������{����������{����=�����{� '.��8?C�{MWa�eoy|�����{����������{����������,���{"(.�4:@D��HLR{�X^d��lt|�{���ｗ��������{����9}��")6=��BEJ{�W^e��ry��{���｛��������{���н�����{������� %*�{/;G�S_kw�����{����������{���������#�{.4:�EPV\��grx{����������{�������������{��!'15��?IS{�Wak��u��{���ｫ��������{����=��h��#{�-1;��DMR�{W`i�rux������{����������{�����������{�"+��4=F�{OXa�jot}�����{����������{������������{$�,4<D��LT\{�dlt��|���{���ｬ��������{���������{	�%,��37:{�ADK��RY]�{dkr�y}�������{����������{�������������sx����%+1{�7=C��IOU�{[ag�msy�����{����������{�������������{����=�� �{�!%��)-1{�59=��AEI�{MQU�Y]ad��gjm{ p 
  %-79�N.>sl��%sc1+M@�SDBL6.0!�zSP�kFc+=�%/vw$u�v�.	txROOT.p?��== ��"O/!/gIN�VALID�d��?:igGPi	� . \ _^  $~!#%%&-{}()@'` �7+�(_�s%s�;:L6P�41 \�����DEERASE4�,lu��
c��
���i�!XR�,u�����^[�|�u��摪݊uc��5��_�lu�z1�}��{	��.����z�s
wW���s�k��W�@:\p3�SP�.k-@FP��v���c`C��(�-�\c.� � sq�/QdD�VS��4V
��etғ	fa5�mxw96.6��6u�S�,5o�+c ���i� A��XTRA$DRVsp6�uu5�WV3_ս� <b�.��yz�Y03uf�) �1�^�4a��x' ���ǁ��� x�����{. ���  ��������������.*��x_�(/%3 �*�������f�MS-�[F������ ������upgr�6] ��w3ipl (�~��*��,���������<'�P �y~"b�^N����  �������7�҅������ �L����������0 ���
���
����3%���04<� � ]�z�ɉ�N�� ��? ��������������|�T���c�Ved�������0���������CD ����%S /��� ��������~.S�NR�94�����$"���-���#�����; &]'f3\��Q	���:�����2����6 6ics ����)ܛ%�܍s�J�f�<����I�wC* �o8A������L�	'(��'�Poك��������R���`.�������̃������ ���8�-��˱�`�è��ɻ�З悃�.�Ն������@�����.� �!�����n��E��� ����x���������������W��������)�̇�->&�"�� ����+���� �ц�����9�ݘ����P[���������.�C���  ����~����B������ ����Y���S���l�X��[u̺̔��l��8�8���c��R������ �N��m�����.���=���9�P���I����>������>�Ƌ�e$�.�A ށ�lud ��P�	)s�k%n�  ��"�0���A�10��>����������G����C����8E���L����O�$��#.D�k���ψ��sA7�����RM\����������	�
j��-e�@9?s^�J."P�MƆp0̑������I*Ci�#�8���H&�˛��x�����������L��ء���.��&��� xe ����0��̅�֠�� �s���ۧ������)�������!�����it�R���!����a����S���  �8�����������ސ��;�B������������"4 !8�9��}�ĕ� 
�n����k�  ����������x��Є����9����q� �ĨB�Q�,1 u�ރ������� Je���������Ǌ�k���=y����V�s:���P�`��: ����:������N��1������2ۣ� �� ����;����!����#3<���<<~�4>����; ?�������`�f��8��$h�������(s�t) ��ٹ��*@ �qŁ��!��Ҡ6�u^ ��U���8h���f��y(�2���3��v���@�p������`�M����'�I*it� }���,��\�������+�4`g�(�e��"�~��-�G��pad �!A����В�M�H�a��a����y�֯�F|N��di���P���de��� ���!e�ܬ��8圐����|`�S�����2�F�Z�{p&;�ă��
 ���ȃ�v��� �0����������)��;����Ǉ����cܘS*�Fix x�'�����WX���b��:t���53^dc����l�����q����Mx �&���Ӏ�����������Dq�ACrAl�&�c�A8�ы�Pp��ǂ������givW̅�!��@;;ꂤ��7���	��2�K�$l`�>���ƈ  ��������form �z�.��(^=,�0~D#�E)N.���5t`�nh��ʽ��ȅI��m<J>�E� =������~pI�la�dU���  ��������������.���#Signa$������2��! ����%ғ��8d��(���9|=Copi�p�upde�{vӄ��M�
�|��P����M�t0Bad � ��a����)ޅ0㧃֜�
"f����6��  `딧����|�1��s�jV�����=�^�y�������o���r���k��`!���� <T8>\:⇍��b- ��*���� �����Ǖnewer ���ÕpT��n+�y �iou�����T����S�����appli&X �fua yirU<p�����XUnAlX��� x������򈂐�Q���e�*d"R dATIO=3 %1:  +�������.�������=��� ��������)9�'�u|�A��2G�􊎫{�D[��'�Ï�"����!�� N ���Μu�a,Q��x�w��6�� �*��#q�o�E������D��������;&��8����P���a� 0Յ����&� ������ρ���q�W2�J�jӎS�k�J�  �PC-��������� ί-���softw04*�Stop ��큽�)�b,O�m�(��ߒ|���I�K�$�SV�Cl�?u�ኅ�����������eAt ��ҥO��#�jB�����%N��2�� Nrtroy ސ� �O���晰���Q��Qh�����������B���sm l����ј߰th�N�p��p�causQ:  m`�-��՘�D�ه�3�U������;�t���N��i �/�a� Ii$���0�����?l l����o�������~���!�
�י��4����~�����<�S%1 ���D:u�K�5����
�R����\+��8��Ï��摏X��X��A�1���A��M�B������/�$�g/� �0�P��]���Ɔ�NU��gM��0��+������{��@Y��Qt�0S̤����Ƙ����������SI����. �E�7��$$�2�ӫ@�6�0`x8����������p7���$��Cx}��Occa u4�� {�������we�K��c�2��@��������+�:�gathe'N�x
��|Q�.��
]��š],���wTt&�_i���2B�ZL���+�
*�!�����ѧ�	����ޕ����n ��v��������������U윻��f�]bw�R��Eg�bet�e n 512 �819�ۈ*������Ǆ���P����.��mark F�����{�����Pi�ㅆ��Lik��p�݆�֜~��;� �������3%Â���y��ǈ �5�Ǜ)0���c����#�xp�y��8�)�� �ek ԯPTC���LH<6`������!-���m��d������hP����Y�$�3��'�n�/��킐���"�J����o����E!��©㍝2'A � stoڕ�w���� `����T��J�����ƕ)������uR.) #��F��Ѳ���K�#ev x�though �d�Ʋ����.K�/ޜ��R��lA����V0�����*�:����6.c���=�v����Q�Є�!�R���LR�&c�q�Cs���;������c���L�����'�; �$e*!�"�8��SFe�����b!R�ʅ-�������8�ˏ��)larg(����+�rand�(om �5d�e�min���"�S{<��W���\����0�޼?�TP,�8I	0w� ��#��H't !�M�U	f
}�0���navi����B�eaddi&��ч#²���2	�dr%Z!�8�z�
��beyt$����c�  �o ����ߒ��88��؊���g�$��Any �ᔧ�5�����������+�
; ����� ��/�������a�������AB�Ѷ�\�I\�����!�N1.��3�}���:��oF�����C"9���U!|����8�+�Ren
IX��ӂɩ�e�ȭu�������1s�*����'�˓�0UŔ ����G�� �����!ҁDIRn �����������������������J���A!��JPAZ �lim���z�2�Ys�����ڂh�����㈊R��!��F.K��6�M%��s��.��
B���-[�!Y��إ�^�tU��i7~��#daB����ul+�`|�������ߜ �ၡ�oT�0����='�6�,�'7J����f��fai�r�	��m�����n��&��eK��g�N�on.֥�>G��B&f�T��t�#�����'����ˉB�5*��E*L%�+pP���>�ܰ��=�Ͱ�����$u}th>	is��D@�
m��(�Zl��%�� ��t����(fW#)�$�������u��n�CB����[&:�b�q��	p�)����ꑩ��� ����&�������*�n�쿗ѐ>�qN����!�yY  nNqQ�j�Oq:=�CRV�U 2��
ou��Sp&riv� C=SCAND@ISK.LOGN�UO.DAT"�qINI(m���)  �b0]��h���.
�C��7!�Q%% ���& i�`�?��z�2��V.A(q�(������[ypa� �|��!�/�3� �%In��׮
ұp�Vd ��������J��||�`<������/un; ������f	�]J�  ���0ܔ�������r�N�9E���$�ޫ@��l���:
��`
�nr��� �
�������c��4:�wvjt�7 �I:%M%p �%�A��B %�����It�c:u���TOK8�R Y�No����P$�rev�S�|en �����4F����:O��o�
"�j�AB���x�r/\ PD ,�Nex>{��"�All{�y$0u2 ��	6	� D�q�lView \��Sh  OS/�Wi��lw�Fa>W�p�@N��@^@�1bcke�Su#�r�r�A�Disk$XtraU�<x��<�<��Kڽ�
�
�c	�(Jip��^d2��m�����3�3�	���	�	�*�	1	��		��	�J��	%��	*	/�3/
" 4
	"�;	�"�0�s	
=H	��T	V	�=����>U�u����^<v ��e�xa�����baA|\ ���  $2 unS�� ��
�0� AW�I�W�;���ai	2	�3�W	>	�	O��	]2-w2TU-|	�UU�ԥ�	3	3TU$BIUU	��UU��U��	+4�TT4YU��)�	�;/����&�R&�	5R�5��	5j��o	���	�$ݪR�	6R�?6D6I��w�>P��	�	��<	7	6	���;9	O��Rr��u����	��T)\�	8U�	E	o()	�8J�8UUn��U���T���8�?9%�{�A�/�KyZ9hT*x�T���T���N:S:��[����ҪI�;I]";RUS[�US��U��<��<>��Tz���	S*	�<��<zU.�U��	=��% &#=�zA	�zU&�]S�Uz�>��>$ݫ	6��J	i*U% &��w�>�UU��	�]�B�0r⎅��x������DӪ�=�	?�t	O	�?���8��B� �|F�2� z�ο�A�JI	@	m@S�TJU�@T�	���@z��T�B	/A�B�ʕ���.9&������ݘ��������as���֕���ݥ�O�*�+�ܵ����ǥ���K�S~pJUXApd	]E�y z���z��S�K~uXR �v���ҡɓ�ÏfK�p.b�JIY B	KB�Cb����u�`�����z2�����nK�O�g�z#��և`�R)~zUUu�	�O8~��ͻ��[����ڛ���~$�a��Y�ݪ�6�MC��	7	tC��_�՘�r�O�0K��_�������]���1��F��<n*��:�ݦ��\U��~�U�	�	D��	sDn���������p".C�(����*�ӂ�܄���ER���0NM�%�;"h�) ��F���t�ؼ�nBkr�ers�oGpwG�ט0���[<����-2�&����1��
����
���F�����o?��<�+?P
ӏ7
7��&��&
vaw�lHčst
��䪀�ER�		dE.h��Nېto�ݲ�N�����;_��toH&�d �mr��H�U�������d�	�+�m '.'�)�0�6q�u]���M�O������s�� e��FT�[	KF�l	蔇��^���!)-0��J�0���x�ωw�o1������
��i:�.�� �XZ�F�U�	�	G.)U.@GY��	�GTU�����	H(�Z-HA�J	t	�H����zX����o��@���U�H�	I^�d���or ��E����B@I��9H	u�	�K�����C
	��� �М����a��MU�b�PUݮ	������ ���������nmp?̣j�a �׶�����aܔ��v�y�f'n<affom�<b���� �$�w�O�(* G�T������B���; hq3Lߍ�s�^�R��ِ�Μ��y��8��T��3����12t�� ���ο�Ի�j���c�|���.�R���������p�%ҏ����'g�Inw=cԐoܞccuDZ������B�>�k�S2ӹ[ˋ*ј���B����&w��C������Oo�]S��t��d딲�nu H$��邗��be��#����+�?�n���8��^c�5������"����{s; O1��'�,�����Y�0�����wde݈a���4� [�؉�јX�(�j�p��������:��
��X�����\�U�{q[����ӻ��F�/����C�0��v����z�݆�O���*|ݦ�y����� ���especiy�o�pq���T�eq/)� ������޼]l�������;���������ә������w)�04���n����ɉ���r��B��r"��Ř��0aǂ���'�V釕@v�'�"��w���>o?g]��#�ܡ����c�+�@�v���ܝ���/8 �k���� �"���\����y�������݆����`�������v�
�Ecv�� �w���������ͱ�l��/8��{��a�ʍ"A C��x����� g��X��������P�z{�	l��?�����ASo����ȀW���fromN@s�����0��?�������tri�E[d ��<N���ac=|R� ,�gene�r+?̋��	���=#`9ma��V�?��$� �����w��L!޲���c�4�q� �|�L�	%��a�ys9��a�ppPnt 5��%3, ��p۷����a� 2������$0p��D����������-� ������v���#X�����f� ��A�futui���c����i�[mprov��yncAe���9��f+qu6A���� �������x������#S����NK������ �4����ݵa#��������d�M�2+��L8�׵����t�~���s���C�liab?�������������[�wD��hIe�����@��safeguOƉgR��12s(se"�ch(��sRu��p����-� gra ��������ǂ��
��:`�[�  : | /�] [/�1��ODn�]��]�p1��B:�����43w\%S._N~3�p3�i!{��{��`/FRAGMENT,�q7][p�]�����������ND,�% ��, �q��[�F�дmp��j�� B����loc������ە�	������mp��01�0s���:�< ���CUSTOM �p��r(���Aordh��\E��tNOSAVE/�Pp��c��r������90�#UMMARY&�&1�*���a�hpHY�summary s�@L�/�ַP�����������MOQ��J��c�mon�h�e ���s?��˛�� �} ����$��E.����r�a#��}tiN��y�������Zbr�����F��#�����afyz �g�s�quick`��K�	|A logi8�talr�`��!�e�Exp��Ms� S��{ce:0m�� �%3 P��%5X�1$~6�ԝp��cT��{�d AT suppor@(7�Õ��w�@zu����ҕ�� �(A��K�f��D��Ɔ������О����< ���(����2��%.��@�{烝��ݥ%S�����`c��3ǆ�mAܓ#��R��%N�Rz���<�1 �;�����%Қ���åi.Ƃ9�)��+�c"��q,�|��
��_��9߰� �O��8`¥�����d*a.;��x�8�lg٫��Ta:� ���j? What ���wh �x���first?�: h���Nn=>PH��� &��s(��CVFsB�{��urx` ���ib�������9A��������^
8t aCheck0����en�	堁 ���X���2�����/0��,Hw��.�lxs�%�
�N�pM���)��r���/��;&�Յ/|�F/�.���{cȀ�MΪ����~��m{����*�*�b}"�m�h��igh�h�.���o��h���D��ͻ���L�"���xyh�� ���ՠ���u���a�����.[�Ϊ'���<��X�+adj_��<��:���?���qUЈU� �>�M��H�� ����������L�e���$�/���#�D�"����������;;[���"M�H��u����:���������晪faP��90;-IfR���&�d%;�t�d3���� 8n�%S /���!��ߍ�#� ������(ά��nCp�'~�S��5Ej��\��un�W���c 	�cE[��'�-����b�����Dh}x���r������
߰�������<�����t��.ǂ�u��t�clud�#��Y��	����:=Fʝ�d�������q��� LoT�ԅÌ�<�v�� v���� , %1�s�U�ρi}(o�	���`��D�xR�����^��oLO� %�Ⴔ��.Ä�����V����#��A	���{�-�����0]e��Å͸	-`�� <��?��Ξ(���)�� YA �B�o̳����� butt�J���H�/E���<�w4��c��l�b��C6{������!S����,�l"�������[���� T~nge Y�y��������Z����2���r��S��B&N}�hHTA��A|������l3��$��Ȝ�pair��]g"�3.�d����b�p��Ģ	���p=Bmak2����@�!���CL��.������  �$b�����������Gfib�t C���ތE�[�Ť#�fy�K\x�5�x��CP�m9$�L$ A:)tP���r5)j�EI�i����_��lg !����Z�*����D�����ʇ�������!��yDX ����'�~���la΁be)!����%]��,,� ����� �IMPORTp�ANT: \����8p������in�2��<U���Mst.�����7��� FQCau�B�ϴ���H��l����eՓ<@�^��)| O	�Ċorpe�7������b����#<a_�a��61A�ۊ�����\f��b��K�ۧ���.�;��k��p�l�����S� xQ��#�j�	@�a�7���=����$��i"�������T��[��]\+lD\	Tmk\	J�8q\8{Jo	�\�S����0�����gWY�X�ӣ�;P�%҉d8y ��ms�ax�S��=��r��GuK*2AK����˔H�R���]��	M	v	bUƜU��	^�9	2	�� Ƒ������������%���e���ł�C�Ү��8 ܾ��������6�4������t2���&�3fX^�*fy	�}l^����_��	I_&v���	�Jo	�_;�`���	DJo	f`���v`"��*	�	�]`f�.�ʻ\٘S;$����I�~�.C��*�V��a	G	r*]	�a��l���v���]��������@��#7����΀�t;s ���y �should�WD܆���������Z.ev�����N�$�A�H٥����
��QUJǝϥ�	b<榕�M����^>lӣ���&mL���Q�o[�_���D� �����]to ���\��������� ���1�\nOAfp ��Q���s���1);���~��;�\��F���i�$^+$tpidW�ߕpow�����
�̔gn 7^�+�09�>���BackbnД������1 S Ȣ��ba+�+aH��rvZU��/�Gug>T\���d\y ��wh't	;7J/�6���ϊ���ŕ��Difi����y�chniV�in�NP���O���s�����]����-���{���䆹�-����:��$ژ!�&bЛ!b��B3<�y	2wT��2���S6�W� l8�ė���܁��/ ��!���+��: �	�	�WU	�	��T	c	"UU	2	L�#	^	 in�	Q	����	���	�	���	d	S��	l	�	���	�HELP*��`
UNDOCCKO`�NLY �p��6`� �������1ITI: �􂏲�������(s) �_��Uou`��ּ�0nMn b��k�����itself
< ��U�
�	�E*	�	�<���_��d*���"zAͤ'�V��9���Di�unnae)�\�-(�0ݝB �o 	=& en�7wz2	�	,e"�D>eDT��W�	��{ B4�������n�*ex����_����N��؁�x�u�0�h�>��_>���: Yo$�齈x�\ �@�/�����i��N`c.����`*�.�L.�t=�� ���3nd��E�na���v'@�Is�R��@�B���� W7���q���5����(�ج
0� �* �? w���dcQsY��E鸒å��|I\C�U/��{��(� X(MOUNT=%3 %2��1��|��8A
�mb-�����5�sx�m��<#�ex�siҘS+� ۧ�M���both�N{��������������� ĂJOIN�������͘�95d���^�������c��-%(�����&���'�������%�VQ�������+UTERLNK��[etwork =���%��Gn�`��.�a��a� �� "Z��� �L�?�=: /%s7�I�� �����$�� ���8�쩉�4�`�{x�&��O�
����

ne� ���F-­ ����r��2 ~Ar� L0���v���LE�,����P腠�����M� ��}���P�I�sp�	��fu�	�R��j͇�)�room ���]�f��A+e���J�"��@.�%y�#�p+�In�ۢ �eNV	�4 �A ���<���#���7x�}vŹ��M݁�*c�����2��3b=�\�4g���/��`bunmod�t ���Due�� �7�9�2�� �h���!�����[�������f��"shed�O��s�(%�x����+ �������rha��������Rp�2 ؏ ����!0�xdeep�ex�=Õ���A��6�����ng�����֥�&�&�9&L�©�cU@#��#H	@"���������ءu����ֆ�����^'z�}�Y���x8��n��8?�O��g�p�� �ε��jϑ�Eu�z儉���>�ѓ���� 4��������Ք�unav��� ����ц��DRV  SPACE.MR1 �DBL�[BIN �ʈ�%x$2.

S���@�����㯕����6ep�"�je��te���������
�/��,I���$�T�����I��we(���e��
ifR�r*	`f.1�TBmfB�U�	�	0g��T	BngT�Kx	�gk�T&����	���&ʺ��T���ggh�.	4h��p

9Oh�wB[hBUUv9�	U��	 iT��iJ}ҵ	�i���X�|x�F �8�
�:
�
U�j

��
@

s Iv�HB��V.�����t2O�����] ��O����& � �fld� �Ro VJM���	VV�RWdN��f���:
����}����,��\ ���­���*�������1�y<=���'�b�v�,�|�,��c��"�d����� ����
�"��
���˫� �G��(r�����&��KE}P@`)#���A���=R�ej
ij6�
�)lg \��Ă��fults: ߭��z��3� ��8� B͎����gr3`��� ����IFF������
� �B����e���6�ގm�p���y��1�# �~ld-�$�r�s8��΂��N�D�c��rZ����6���
��z��H(��.��`�V�b��%1�&T��䤂��(�Y7
nI_c�}�D���#�2Ꙙ����Z�V|��#rB�i�a�dY�8�t��+�e�|�o�p"�����]��Sǥ~;it2�� �˔�n�crT��k�:\���Tr�̯���h�ꠑ��| ߭۟��X߹2��XGW���~t� �>������
������DOZ��3���;)�������v�Z?����\ �bj�(�P���2<����R��.�%1 �����\A&��%���74�[��~��qZs�tګ�����>T�T������0N�z�^�^����CG��:ݢ�o��"��]���=�2 dout��������M�n�"�ʁ��patch@-֑HG�.M�J[���.Vx/Ã�~;���xU�	�	���	�;�)�������W���r7�0�W߲��͞�s=�)���K-��� 	K<v�ꊢ
�
	r�U
	i�)�	k	A	:�{ C܁�@��!�(�YkL��|	�k.1UU`�N��}	/lW�R&HlKU�	�&�k��J'��p.�޴�KX���������NO���ve(o�~ n�{�mad���q����յ;�,o��̦�3�˪t��	m���)�tP=�܅��ձ>�����~�C<���S���V2�'6�Tm�%Rj	M��:~	]S��� �mj�*nV	O]Cn&�N����{����; @ۓ������{u�n@9k�' �ENVIRON�Ó�0~AUTp�OLOR DELET3�rFIX3�OFFN�fP1MP�<QUISAV$SK7�I�NE�8ALWAYSLPP��WD8WR,�N'D�n4 Miep Y8canTimeOut �L�Chec�Pk�fn3
NumPas/s,�urfac8Ho��s2Dr��hTr��UpllSa�� �RSp6Rp���ff�6S_Hecr ���e_M�aƤk�_���_n�_����Boot_S�Uo,In��vZd_�� �QBGt�S�\�^u}���mS'e��L0��>s�^/ %c:\�$ 	TH]= C"Oz�S\MS��6_Zs\ mrc�!i.txDWA.pܸ=== 饸y B \X.XD�PEC 
 	#;[]=	�^�d ��_FIL�E_sFO= � � �V �"%�p�v�14i��� ���� �؋�*� (� H����T�_s ���F h g��Sun� Tue WedhuS��iNo�t��Cy("|�
(s�_.n4r��:(/e@Ja�^FebDar Ap�gJvl�ugfp ODcnNov Dec0�Eu56��r<ch>��Bil
M�_iNeU�
l��Z���`temb`E1fo l�%r
A M P܍u2\ 6+0&�&��%�g5�/ 9	@���XS��
&�E50e�!  0PX< 0SWP8�S`yޛpx" ��(n�<,)_D�{�"}�Q.�TZ0#*STD�p��ȏ�̇����p��8������xq�pjc8\U�NG@ |� e+�	`b010203040��607080912X�M61�l��p� ; � � � � � 0ND m: Y w �   � � � /Ml1��#SNANQ�R��D�Nk_`�2 �f$�7y�ACH����Cɥ�E�	l�-��Ȓ*i�/�J��61�/�<u2V{m��Z:.�{{�4R�f$r��F�^�J{�
�kP���l'�J��ҽ�?�{F��l�?�C�^��$�d����~��v���
-
ƽ<<NMSG>>
R6	܎
- �Sck �pIrflowM*&3��q div>x by 3R 	!9!not eughHٽ� ?�Q.ronm��>.�č�� ���-��v�r$1�AE2Ex�ng��-poq ��\�K6A��/1tN�+���_�\k� : M�k�U:�v e i�s/f �}�{�g ��h ��i ��NjD�ѳcskem�0=ul�� sq�F�(�m��n ��do�pWp�xp�cit���g�<�U8  ��; 
  *  �������j��������|uV=,'"� � � � � � � l d [ V Q E . )    �;          ��A�������wpg`�;& $ "    X| ��� � � � � � W < # _G@3,
���pi���md]> ��mf�
�
_
X
�	�	�	�	�	�	r	a	I	+		�������\>������uL�zpf\TLD<2(�;D B @ > < : 8 6 4 2 0 . , * ( J� �;H F 
J�o;���r\L*�;J 4J��}aT'	�
�
�
p
f
J



�	�	�	�	�	g	I	6		 	�����qg��wdP7����xUC$���;L Jvo^JC#���tA&��aMF/ ����;P N )J���aSG����XJ>����K=1����F����YNB����{b6�;l j h f d b ` ^ \ Z X V T R &J�0��j�o�K8wP��gF��O(!����e^PB4&���;n J�!s!d!U!F!/! !� � s D  ���Y�;p J�!�;r kt / �;t v k,�;x z kJ���;| koX�;~ k8�;� k��x�;� kS7,����{tUB;� �;� �@����aJC���	�	����.�;� !�vKD/ ��zC ����
_
�	�sbV=, @.�������;� 	��Y!��Q���;� � � � ��}o_-����_5� � � � ( �;� � � � �M��;� ��cM	L��
�
3

 
�	�	t	P	I	��s�T�;� 
�� � � � � | t ` U / �;� � ��;� � ��vnT�;� �;.%���
�;� � � � � � � � � � L�����tG�������O81)���i�		v	n	f	^	T	L	D	2	'		����������sh`XNF3(���~vME����yq80�;

�	�;� ��
Z
�;� � �  �/ ��������xjN)���fRF:.��HA9+�
�;� <����yG����a=������h]RJB6+#�X���uhJ?.&��������qJ������j-	�;� �7*���;� � � � � � ����;� *����{cZ<5$���������m9����zs����������;� � 
����tP:)!���;� � � �zpg2(��;� � � >���5���$�"�"�"�"I"""�!�!�!!	!� � � � � t < / ��nQ&B&/&&�%�%�%�%^%R%4%�$�$�$�$`$$�#�#�##H#<#0#$### #�;� C��*�*�*�*�*�*]*I*&*	**�)�)�)�)�)�)�)�)�)�)�)^)S)B):)2))))�(�(�(�(g(9(((�'�'�'I'Q.8.�-�-x-G-�,�,�,5,�+�+q+O+++�*�*�*�/�//
/�.�.�;� � 	��0y0l0d0P0H0/0"00y2���������zvfbWRC>:/*&���;� �����ZK2���haYF*� � e B (  �;� � �����mO���kA+�����;� � � ����zTM0�;� � )��	v	j	O	C	&	�������p^,%���~aD��������G3	
�	�	�	�	�;� � =��#����~S��J�
�
�
�
s
a
/
`;.'�����t[S(���iB�����>,�����tb?������; � �	����� { [  �;�	qW��XQF6/����;
�	w$��m^2��cH/�;#�	�
�
�
r
\
*

�	�	�	�	h		�����]@#���~W����vL2�;�	��RC��������xb1*"�;$�	��hOD"����wphX-������xQ�����R ����;�	���gC�;"�	 >��oY81)�ykW�A��!i >  ����>�;�	�$�$�$m$K$$$�#�#�#V##�"�"x":"""�!X!�;�	]%C%%�$�$�;#�	)�(�(�(:($(�''�&�&[&A&$&�%�+~+c+I+/+++�*�*�*�*n*G**�)�)�)�)�)q)M)�;" 7�	X/,//�.�.�.t.>.�-�-�-z-i-C-7-(--�,�,�,~,',3�2X22�1�1S1311�0u0h0J00�/�5�5�5d5<5555�4�4�4M4(4�3�3�3|3W3;3�;(&$S&��zg&�;*SEL_�;.,0S 	�;2Si
�;4S�;6S��;NLJHFDB@><:8+���� �� � � ��;TRP+���tmb�;V�+9��>%��}N5+����k?�����5������e[5"������x]J.�����lP4�@2 ���rCwfK��|ZD������vX"0""�!�!�!�!�!h!K!#!
!� � � � � � � v Z I ��/_&K&�%�%c%�$�$V$�#�#=#�"*�)�(�(.(�'�'�'�'w'T'�&�&�-�-�-�-w-�,_,=,#,,�+�*g*E***1�0?0�.�.�.v.�-+22�1�;ZX+t4h4/44i3�2�2�2�2}2^2W2r� ��;\r�v,���
Z��kX��=��Q�y2���|xtplhd`\XTPLHD@<840,($  ��������������������������������|xtplhd`\XTPLHD@<840,($  ��������������������������������|xtplhd`\XTPLHD@<8�!�!�!�!�!�!�!�!�!�!�!�!�!�!�!�!�!�!�!�!�!�!�!�!|!x!t!p!l!h!d!`!\!X!T!P!L!H!D!@!<!8!4!0!,!(!$! !!!!!!!! !� � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � | x t p l h d ` \ X T P L H D @ < 8 �y24 0 , ( $            �����������������������������0$,$($$$ $$$$$$$$ $�#�#�#�#�#�#�#�#�#�#�#�#�#�#�#�#�#�#�#�#�#�#�#�#�#�#�#�#�#�#�#�#|#x#t#p#l#h#d#`#\#X#T#P#L#H#D#@#<#8#4#0#,#(#$# ######## #�"�"�"�"�"�"�"�"�"�"�"�"�"�"�"�"�"�"�"�"�"�"�"�"�"�"�"�"�"�"�"�"|"x"t"p"l"h"d"`"\"X"T"P"L"H"D"@"<"8"4"0","("$" """""""" "�!�!�!�!�!�!�!�!�&�&|&x&t&p&l&h&d&`&\&X&T&P&L&H&D&@&<&8&4&0&,&(&$& &&&&&&&& &�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�y2�%�%�%|%x%t%p%l%h%d%`%\%X%T%P%L%H%D%@%<%8%4%0%,%(%$% %%%%%%%% %�$�$�$�$�$�$�$�$�$�$�$�$�$�$�$�$�$�$�$�$�$�$�$�$�$�$�$�$�$�$�$�$|$x$t$p$l$h$d$`$\$X$T$P$L$H$D$@$<$8$4$�(�(�(�(�(�(�(�(�(�(�(�(�(�(�(�(�(�(�(�(�(�(�(|(x(t(p(l(h(d(`(\(X(T(P(L(H(D(@(<(8(4(0(,((($( (((((((( (�'�'�'�'�'�'�'�'�'�'�'�'�'�'�'�'�'�'�'�'�'�'�'�'�'�'�'�'�'�'�'�'|'x't'p'l'h'd'`'\'X'T'P'L'H'D'@'<'8'4'0','('$' '''''''' '�&�&�&�&�&�&�&�&�&�&�&�&�&�&�&�&�&�&�&�&�&�&�&�&�&�&�&�&�&�&�)�)�)�)�)�)�)�)�)�)�)�)�)�)�)�)�)|)x)t)&y2p)l)h)d)`)\)X)T)P)L)H)D)@)<)8)4)0),)()$) )))))))) )�(�(�(�(�(�(�(�(�(�;`^3i��c>0!�����xYD2������rkD� � � p i R : / ���1��=-#���;jiX	Q	�����cP�>I1�
&
�;li#������;pn*i�A��Y���7�nS��>��za�a&����e[K�\J+�����}R�;ri=(!������~r^F:�;vt?I�=![� � � � _ A �;~|zx?1�$��;�?-

�	_	(	!		�������
b
[
F
�;�?c*���;4��*#���+����;�*?Y6��e^I!����~a0$����WP0���xG��l!�VO
~$���0���{X?� � � � � | h - ! �;�����lB�;���j?8�;���p/!��jJ�����;��	���H����c\4-�;����R@��eG�
�
R

�	�	{	�;�����(!����9��o83$�;�y2+�;������� �xm\S5����xmP&����ypR!� � � � � � j @ - �;���k9��;�����2�			������w[M7��������cMB:*�����bWJA0( �������Q	J	�;�X��������yg9.
����vc\G�
�
�
�
�
�
m
b
Q
>
7
#
�	�	�	�	�	�	��k`YB.#�������QJB)������shWD=-������sE:)�;�B�aYQ�����yngP)��������wd\T:����Q@5(�����ZD7����vYQI������;��������m>6.�����~����������;��������a3�;���VM8&	�����z0�����]	������uK"D""�!�!�!�!�!�!�!�!�!!w!d!6!-!!	!� � � � � � � l ^ V ���PF9,������%�%�%�%�%�%x%q%i%Q%J%B%5%,%%%%%�$�$�$�$�$�$�$s$Q$8$-$$$�#�#�#�#�#�#�#�#�#�#�#~#c#\#P#I#A####�"�"�"l"�)�)�)y)))�(�(�(�(�(�(�(�(�(q(Z(I(A(%((�'�'�'�'�'w'p'/'$'''�&�&�&�&�&�&�&�&�&y&q&d&[&T&L&1&*&&&&Z-O->-+-$---�,�,�,�,�,,h,P,,�+�+�+�+~+v+Z+P+F+�*�*�*�*�*�*�*u*R*)***�)�)1	1�0�0�0�0�0�0�0�0W0E0:0/0"000�/�/�/�/�/�/�/�/n/4/#////�.�.�.�.F�u.n.J.?.2.)...�-�-�-�-�-�4�4�4s4j4Y4F474"444 4�3�3�3�3�3�3r3W353�2�2�2�2�2�2�2t2X2M2<242,2�1�1�1�1�1�1�1�1q1^1O181+1"1
6�5|5s5l5d5W5K5D5�;�^kdSD70� � � r T > �;�^6L�I �;����� � � � � � | �;�������
�����s���Q!�;�������UE9�;�����(��H+�����:�;����
���
�
E
w	5	��&�;�������iV?,��zs]V9��/��{Sc�; �n!��!���������!�mf��_L=�H���;�xW=#���@4��th5%��%!!� � � p D  �;
�w"Z"�!�!�!I!B!�;d�1&$&&�%�%�%�%�%�%�%}%i%Y%L%:%%%�$�$�$�$�$�$�$$r$b$B$2$%$$�#r#Z#9# ###�"�"�"�"�"�"�)�)T)9))L(1(((�'�'�'�'�'y&l&U&A&�-�-8--�,],N,B,�+�+�+�+c+)++�*�*v*6**�)�/�/�/q/[/:///�.�.�.�.{.f.>.7.0.�;��������zfZM9� � � � � v ^ E "  �Z+�;�Ng s: ���q[�;$��B4�
�
�
�
j
R
:
"
	
�	�	�	^	����x�����6J0�
* # �;
� 9 �; 
�#�;"$&
	���;,*((��xiM6������}cO �����~]O
� � � o K @ �����;.6������veYD1����viL6����pQE4(�������;	�����N@2	����;20	��	�	�	u	g	V	N	;	4	�;864?��}eLA6) �����������tc[SD7!�
�
�
�
�
0

	������W4(�����~qP�������;<:5��hOH.������������r;	��~V<1��x\>+����saB(���r]=6
��y2hL_L�L�L�L�LMM�L�L~MuMlMcMZMQMHM?MNN�M�M�M�M�M�M�M�M�M�M�MCO:O1O(OOOOO�N�N�N�N�N�N�N�N�N�N�N�N�N�N}NtNkN]PTPKPBP9P0P'PPPPP�O�O�O�O�O�O�O�O�O�O�O�O�O{OrOiO`OWO�P�P�P�P�P�P�P�P�P�P�PzPqP�PQQ"QQ6Q-QJQAQ^QUQrQiQ�Q}Q�Q�Q�Q�Q�Q�Q�Q�Q�Q�Q�Q�QR	RKRBR9R&RRqRhR_R�R�R�R�R�R�R�R�R�R-S$SSS�R�S|SsSjSaS�S�S�S�S�S�S�S�S�STT�T�T�T�T�T�TuUlUcU�U�U�U�UmVdV[VRVIV�W�W�WwW�W�W�WcXZXQX3Y*Y!YYY�X�XYYPYGY�YYvYmY�Y�Y�Y$ZZZ	Z}ZtZkZ�n~nunbnYnFn=n(ooooNoEo<o3o�o�o�o�o�o�o�pypppgpTpKpBp9p&pppp�p�p�p�p�pny2�q�q�q�s�s{shs_s�s�t�t~tutltctZtQtHt?t6t-t$ttt	t t�s�s�s?u6u-u�u�u�u�uM}D};}(}}�|�|�}�}�}|}s}j}a}�}�}�}	~ ~�}�}�}y~p~g~T~K~B~9~&~~�~�~�~�~�~�~�~B9VM^�U�w�n�e�#�������ׅͅÅI�@�7�o�f�]�����熃�z�q�������هЇǇ�;DB@>Q!�g���}_E4	I �;LJHF
Q!����t7���6�;NQ!]8���k�����U�B�;TRP��!*�3#��yP� � � { b R , �����gL$�E�����<�xfWL:+ ���������{p]NC*���������zk`N?4"���������rcXF7, �����������~odRC8&���������vg\J;0���������n_TB3(��������t/x 
$�������; 0& � � � � �*  y2��0&.��y2������0&a@#4�zv\9�y2��0&���m\H/�P+���; 
  0&�y2��������ĎȎ�; 0&�y2V�Z�^�b�f�j�0&""�!�!�!�!� � � #�"�"�"e"N"y2����0&�$�$�$�$Y$*$�*e o � � =d��0&'*u)E)((�'�''�&�&�+�+�*{*�+�+�+�+	,,S0�; 	0&x0i11�1#33�3w4�8 |<`$0& ,9

LASTDRIVE=Z
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       MZ�      � ��R�    s                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            ���	6�6���`�$ r6�6���k	Ð��]	&�E3�tW&��t@u�0�u�?_�?	Ð��1	6�>+�+���+	Ð��	6�>���6�<�~�	Ð��	�T�\��*�V��� r)�6�>�6��&�=u����/^V*��s��^������.� ��u��� �V r��s�! ��.� ������L�D�t����.� ��u&�}3 t��� ��s�! �c����H �U&�}3 t5W�} ]r.�/r$�m
�E�E�]�M�U�D��|6�<�E��	�$ ��! �]�&�}3 t3W�7 ]s,u*�59l
u#��9lu6�.<9lu��.�  �.�6  ���s�! Ëڒ����t$��s���u���� V&�u3V� �^]�3�F�! �����WQ&�}3 t,&�u3�D��t���s6��6����+���+����! Y_�VÐ��H�\�L�����
�< t|$�It��WV����
�u�^���|�I�}+�u�_� ��ËE���t+��t;|
u;TuA�4��ڋ]/_���Ã|3 u<6�>�D/6�<�D1�r(�\3�L�����;�u;�t�w�W�ډ|+�D-����P��	�"�
�< |t���f�|�t�&;E/u
&�M1#�;�t&�}+��&� PSRV&�u+�u^t�< t�V+�6�>�6��&�E-V�5��/_^Z[X�u����&�u3�\�7�t7;|
u,��;Du%6�>:]u	6�<;Du��.�  �.�6  ���ˋދ4�������������������������������k ����t���A ��.����w�t+�K �����
�u	&�m/;l/t� @@������r�t+�ո  ���Ê���$�<pu2������������*�ËD� �t��������pu$ �����t��Dt�� �V��
�t +�*۬؀� B"�u��
�< |!t:\tt���_WV���^u�XX����"�u^�� Ã��
�< |Wtt��D;�s���+�= rS���  �@+�[ЉT�\�+��������.� .� ��ʃ���^���Ë�RS� [Zs�XX�$ ��P�
���L�< |=u;�tM���;�u����ߌ؎��W��t�]3�}+��_� �u)}뻋�+�[+�Ë�DDu	��� � �P��	�vVS�
�\�< |t���8 u��X\��[^���&�]3�w��t*9|+u9D-t�t+��&�E+�D+&�E-�D-3�&�]3� �P��	�#���|�5#�tb��u*�l6;.<u�t
&�l/6;.>u��6;.�u6;6��5t��+l��lr�l+�l�s���5�3D3\3L3T�����! ]�.�>  #�t	�5.�  ��$ ��VWPSQ6�6�3�S��/[rF��/tC���6�$ � ��C;�u���, �8 ���u��>  Zt�� C����6�0� Y[X_^Ë2 �>4 ��t�&�E������.�_
�&�= t&�]3���;\u�\���&�E�D&�E�D&�]3����\��ÊD$�<puw3�S��/[rl��/t*&�= t$&�E;Du&�E3;D3u&�E/;D/u	&�E1;D1tC���  VWS�>���X_^&�3�P� �/Xr&:tC��6�6������6���PSQRVWU��6�2���rI���w6�<9D1u;6�>9D/u2�D%� =p t=  u"�t+�u׎��w6�6�6���o���/��c�]_^ZY[XÐ�&�]�　t� &�]3�u� �3V.�w�ȸ�/u�t+�tf��v
��u�_ �W�u&�]�\&�]�\�D �t�| �4&�]�\&�]�\�D �t�b �&�]�\��t�|5 u�D  �\5�t+�^� Ë\&�]�\&�]�\&�]�\&�]&�E �t� ��\&�]&�E  &�]5�Q�,�/Y�SV��� ��	� ^[���
�uô���    ��u
�u���.�.?	������������������_�����������������������G�����P���*X�P���*X�ASC: SFT already in use
 RMN: SFT LCK fields not 0
 RSC: SFT not in SFT list
 Share: Internal error
         T	  X	  \	  `	  d	  h	  l	  p	  t	  x	  |	  �	  �	  �	  L
    U
h
  �  
t
/F /L /NC     
t
/?    ��             �
���
�\���F�

�  ��ƃ����  �ʌ�+Ӄ����������V�/5�!�?	�A	�/%�C	�!�R�!&����
�� � �&�>D  uO&�w�|uE� �; ��  ��������&�G  &�W^&w&�_�  ��� ���  &�D  �V&�&�M�}&�  &�E  &�E  ��;���3۹ �>�!C��Z� 1�!�L�!��� r�R�!&�> t��� �, �t���I�!�M�2��/<�u��� �K3��Ë��/���t��� ��&� +�= v� 3����������� ��.�

� ��
�� .
�� ;�wu
;�v��< �	�.��
���.��
 X�м �S��s
��� 3�P�� R   SHARE � 3�3��΀�w&��u".�M.�O0.�P.�K� .;6IvA<u.�M.�KA.�IR���t<	u.�M.�KA.�IR�6GP2��QXs� �H.�>�
uø�L�!ø Y3��!� 3ɶþ� �b�!�۹  �>H
�  &�6I�>=��u� =  u�	 �ځ�
t� &��
&��
��q
u� � L�!��^
u?&�>�
t&��
&9
s&�
�Q� &��
VWQ�R�A ZY_^�&��
 �-��a
u&�>�
t�&��
&9

s&�

���d
t� � �J��<	v�	��.״��� 						�Ȏظ,� �  ��� �  �/=/t@���            ����        ����        ��������    ����       
     
 $A �MS DOS Version 6 (C)Copyright 1981-1994 Microsoft Corp Licensed Material - Property of Microsoft All rights reserved PSRW3Ɏ�3��.� �/.�.�>�.��/.�.�>�.��/.�.�>�.��/.�.�>���.��.�>�.�.�>�H.�.�>�.��/.�%.�>#.�6
.�$.�;  .�=
 �<.�>'� �0 �C Q�R rY_Z[X�����PV� c�!r
.�6/.�1^Xø D�  3��!�����D�!ø D� 3��!���D�!ô0�!=u��= s����� � �  � ����PSQUWR��.�3.�68���t�u�& ��rZ�_�����_Z�r]Y[X�����PSR.�3���u�, ��w s�Y�  �!2�������t;�t� ���rZ[X���u�&��!��� s&�U�!����t	&��!GIu���WPS���ٰ��u+�K��[X_�3��tO�@�׃�u(�!P&��Z Xs��@B�!�&�=u��������UQ����Y�!s�;�t;��u��]ø' � �À��t�ƀu�>6� ����W.�>/�t&�= �t&:r&:Ew�GG��_�.�93ۓ�.�6=�.�6=��	v��7���0RA�u�t<��u�|
,u.�6FA�$��u�|
,u.�6FA���u�|
,u.�6FA�3��3�3�.�69�3��t!�%� &8%u
&8et:�u&��K�sGGBIu�V���t5M.�>; u,�D0&:Eu�<0u�t4��.�>8�uBBIIOO����W+����_Ys�g�Q�ʀ| t�tIIGG�^��u^�	���u3��t>UWQ3�.�>; u�Du�|�q� ���" rY_]^���
�.�>; ur�*�.�;  �3�.�;.�=
 ��X.��?C��@u�
��u�
.��?CC���VS3�3ɀ��u	.��'���(��t	.ļ���= r=' w	.ļ���.ļ��Ã��u���u��.�;���� 3����� t�T ���r�u뚜��u)RUQWP� �/<�Xu	�ظ�/��s_Y���� ]Z�����[^�WP���2����IX_Ã�u!.�>#�t=��uP.�;.�#X�.�#�3ɀ��t&�M�	.85u.�M���s-��t���t&;�.;u�	It�����r����u&}r2�&�G.�5 �3ۀ| u.Ǉ? -CC.Ƈ? C� ]3�3�.�5�D	:�v*����D�t�D
.��?C��@u� ��u�| t8Ls*L�ъL�t%�Du�Dt&�G�X.��?C��@u�C ��u��D�u
�t�D
.��?C��@u�$ ��u��Du�Dt�
�t	.�9��u�� U�QW��3ۍ>?�Q�r_Y�����]�D0u&�PA�8�s&�EP��&�
�tGA��+�U��    4 	 G ,R -� .� /�  =Incorrect DOS version
%1 already installed
%1 installed
EInstalls file-sharing and locking capabilities on your hard disk.

SHARE [/F:space] [/L:locks]

L  /F:space   Allocates file space (in bytes) for file-sharing information.
G  /L:locks   Sets the number of files that can be locked at one time.
+SHARE cannot be installed under DOSSHELL.
�>J����  �� Insufficient memoryExtended Error %1�>���8�   $  / 	 P ��i Too many parametersInvalid switch$Parameter value not in allowed rangeParameter format not correctParse Error %1�>��� �1	� � ��    �     .��  �.��.��  .��  .��  �s���S&�&:s� [�#.�6�SWU��.�� uC��*r<�t7�u.�� u�V�&.��AtN�.�<=u.��C�sŬ.�C�N.�6�.� .��&��6�.�</t6.�<"t.��uT&�G2�.9�s.����CC�&�� �i.�� �`&�G2�@���&�2��tCS&��� [sACC��.�� �4&�G2�@���&�2���@�&�2��tCS&��] [sCC��.�� ]_[.��.��.�6�.��.����P&�� u.��.�< u� u	.�� �P���� X��X���UQ&�O2��t�o	�ws� ����.�.��Y]�&�~  tE��E�.�����rJ.�&��P.��+�.�X.�6�.�< u&.�|�:u	.��	 �&�? t&� u.�� �	� ����
P���� X��W&�.�>�&�&�eP.��&�EX<u
&�U&�M�Z<u&�U�P<t�<t�<u&�U�><u.��@&�E&�]�+&�u&�MP&�Gt��	&�Gt�� X&�Gt� _�.�R P&��uPSRW.��	 ����[�_Z[X���>�� �t.��  �� .�>�	u&� @t.��  �� .�>�	u�  t
.��  ��.�>Ru.�>� u.��	 X�PV.�
�t<:u.�| u.� �	�PsFF��^X�VR��.��=r
�t� .��FF��Z^�<�s<arE<zwA$��=SW�>M��t�>H.8tPQR�e�»��� ����!ZYX.�].�ECC,�&�_[�P.���.�&��.�<+t
<-u.��F� X�PQRV3�3�S.�
�tB�� r92�������� r,�ڋ������� r����� r��� rՃ� � rF�[� [.��t
���҃��� &�w&�< u����t�F&�< t`F.���u&;Lr6w&;Tr.&;Lw(r:&;Tw �2&;L|&;T|&;L
|&;T���	��u�.�� �����&�$�.��	 ����V�^ZYXÜ.��u�Ýp����<0r<9w,0����PSRW&�&�
�u���	.��	 �����_Z[X�PURV�.��rr<�E�.��t<=u&�~ uq�.��t<:u
&�~  u\F�\&:F u
�tRFE�&:F uEF.�E&:F u:FE�.��@t&�G  t&�~  t"&� t<:u	&�~  u�< u&�~ :t��.�6��^Z]Xì�" t�S u.�� t�.��At	N����N���SQ<t-< t)<
t%&�}r3�&�]��&�9 t3�&�	C&:t��<Y[�SQ.�� .�&��< t6<	t2<,t1< u�< u� F:��&�}r3�&�M�t� C&:t��< Y[�.��.��u.�� :���.�;�t
</u����</u.��@��VS.�>� u'PQRWU3��޸ c�!���]_ZYXt).�6�.��.�6�.���< t:r:Dw��FF���[^�  ���& �����=p   
Divide overflow
 You must have the file WINA20.386 in the root of your boot drive
to run Windows in Enhanced Mode
YNyn @M;S<>==?KRRAA   $   (   !     �+��W�� �_���.���� �  � �  �����   ���� �  �� �  �� �  ����NUL      � ' ��� � 	 ���                                              ����E � /�/   �  �  �  � � 	 �� � " ��    ��  
 � 9 �  �  ��   �  ��   � � ��� � , ��� � ] �d � ���� � ��EA�A��EEEIII�����O�OUUY�������AIOU��������������������������������������������������������������������������������������������� ��EA�A��EEEIII�����O�OUUY�������AIOU��������������������������������������������������������������������������������������������  �   ."/\[]:|<>+=;,�  � 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`ABCDEFGHIJKLMNOPQRSTUVWXYZ{|}~CUEAAAACEEEIIIAAEAAOOOUUYOU$$$$$AIOUNN��?����!""�������������������������������������������������S�������������������������������  �<�s�,�S��
�[� �  �Ȧȥȥȥ&   *   )   )% � 3 �l � = �����   � � 	 �NO NAME     &�O � �  ���	
		P 
!
T�VR2	UW	S$&'Z�������� 
!
"2	#$��"� � '� �  ��  "    2    �      �  " �    �         ��!>�  c:\wina20.386     6� �u6�6X�(�>  u7��
    �      #                          ��� .�.b��� .�.f��� .�.j��� .�.n�� .�.r�� .�.v�� .�.z�� .�.~�� �  �.��.���#�y .�.�.��.���$�e .�.��(�[ ��? �.�! �Ћ��V�ڋ���' �!���&���F ��������X[YZ^_]�SP�.�cX[�    �   � ���QVW.�6g.�>k� ��t_^Y��SP��.��.�&��Ȏм��.�c�t.����.�&�X[�˴�<t2���2������<$t	�� ������p      "    2    �      �" p        Q� ��Y�8�  �\COUNTRY.SYS � 4 �� �
  /  �  �  �  &  �  $    , . - :   �  ,; �  �
A20 Hardware Error
$6�66�t萐6�66�t�QW�)��_YQ�<t�.�~.�|�ˎ���3�P6��&;E/X��3�����6�66��״�6�>	�� �t�G��
�t<t��_6�>6�_���<$t�������  ˭ �� ��������    p�;;RB��� �  ��� ��O����P�4 PˌÌ�H�؎�� � ���G����H��� ��������+�s��+�����ڋ������+�s��+�����¬��N���F��$�<�u���<�um�¨t��2� �3ҭ�����Î�������t&��� �t�� �܌�@����&H����Ë> �6
 � - �؎��  ��֋����.�/�@� � �ʎں�!��L�!Packed file is corrupt 



"
&
*
.
2
6
:
>
B
F
K                              ĀtC���R
 �Du�R
 �(&�&�U�Du�ƀtC���R
 �Du�R
 �D@t)PR�82��T�!s�[,�D
��ZX�D
,����ǈD
�����t3Ҳ-RU�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               MZ" "     � ����    �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      STACK   STACK   STACK   STACK   STACK   STACK   STACK   STACK   STACK   STACK   STACK   STACK   STACK   STACK   STACK   STACK   STACK   STACK   STACK   STACK   STACK   STACK   STACK   STACK   STACK   STACK   STACK   STACK   STACK   STACK   STACK   STACK   STACK   STACK   STACK   STACK   STACK   STACK   STACK   STACK   STACK   STACK   STACK   STACK   STACK   STACK   STACK   STACK   STACK   STACK   STACK   STACK   STACK   STACK   STACK   STACK   STACK   STACK   STACK   STACK   STACK   STACK   STACK   STACK               ����        ����        ��������    ����       
     
 $A �MS DOS Version 6 (C)Copyright 1981-1994 Microsoft Corp Licensed Material - Property of Microsoft All rights reserved u � 	 �\ � P �A:\ � P �B:\ � � �\ � 
 �A:\ � Q �A: �? �.??? �  �? �.??? �  �..   A:\ � A �B:\ � Q �B: �  �B:.. �  �                               & � % � � ��PSRW3Ɏ�3��.� �/�
 �> �.��/� �> �.��/�" �>  �.��/� �> �%� �>  � �> �3� �> �.��/�* �>( �; 
�� $�@   �B 
 ��>, � �. �A Q�P rY_Z[X�����PV� c�!r�64 �6 ^Xø D�  3��!�����D�!ø D� 3��!���D�!ô0�!=u��= s����� � �  � ����PWU� r����t���]_X�VS3�3ɀ��u��, ���%��tļ ���= r=' wļ ���ļ  �Ã��u���u���@ ���� 3����� t�T ���r�u럜��u)RUQWP� �/<�Xu	�ظ�/��s_Y���� ]Z�����[^�WP���2����IX_Ã�u�>( �t=��uP�@ �( X��( �3ɀ��t&�M�	.85u.�M���s-��t���t&;�.;u�	It�����r����u&}r2�&�G�:  �PSQUWR��8 �6= ����t#�u�/ ��rZ�_
�t������_Z�r]Y[�������PSR�8 ���u�, ��w s�Y�  �!2�������t;�t� ���rZ[X���u�&��!��� s&�U�!����t	&��!GIu���WPS���ٰ��u+�K��[X_�3��tO�@�׃�u(�!P&��Z Xs��@B�!�&�=u��������UQ����Y�!s�;�t;��u��]ø' � �À��t�ƀu�>; � � ��W�>4 �t&�= �t&:r&:Ew�GG��_Ï> 3ۓ��6B ��6B ��	v��7���0RA�u�t9��u�|
,u�6K A�"��u�|
,u�6K A���u�|
,u�6K A�3��3�3��6> �3��t!�%� &8%u
&8et:�u&��S�sGGBIu�V���t3M�>@  u+�D0&:Eu�<0u�t4��>= �uBBIIOO����W+��
�_Ys��Q�ʀ| t�tIIGG�^��u^�	���u3��tVUWQ3Ƀ>@  u-�Du�|�L��Dt�Dt�Du�|�Z� �R ��  rY_]^���
��>@  ur���@   �3ҡ@ �B 
 ��X��D C��@u�� ��u�
��D CC�� �3ۀ| uǇD  -CCƇD  C� ]3�3҈: �D	:�v*����D�t�D
��D C��@u�| ��u�| t8Ls*L�ъL�t$�Du�Dt&�G�X��D C��@u�A ��u��D�u
�t�D
��D C��@u�# ��u��Du�Dt�
�t�> ��u�� U�QW��3ۍ>D ��r_Y�����]�D0u&�PA�h�s&�EP��&�
�tGA��+�U�]3�3��B  3��D u$&��Du��tC$�B 
 �Du�B 
 �T�Du&&��Du�ĀtC���B 
 �Du�B 
 �(&�&�U�Du�ƀtC���B 
 �Du�B 
 �D@t)PR�82��D �!s�K ,�D
��ZX�D
,����ǈD
�����t3Ҳ-RU�QR���v��$�������!��
�t�e�s�Ȋ��!����� rZY������9 �  �  
  o � � �	 �
 � �  $ 1 C Q a n { � � � � �  # " 2 3 6  :! ;" C# L$ Y% �& �,�-�.(/T0�1�2�314_5�6�7'8^9�:�;<)=k>�?�Incorrect DOS version
Insufficient memory
Invalid parameter
XDoes %1 specify a file name
or directory name on the target
(F = file, D = directory)?&Press any key to begin copying file(s)Path too long
Invalid path
Cannot perform a cyclic copy
Invalid date
Unable to create directory
Invalid drive specification
%Cannot XCOPY from a reserved device
Access denied 
Too many open files
General failure
Sharing violation
Lock violation
Path not found
Insufficient disk space
#File cannot be copied onto itself
Invalid number of parameters
#Cannot XCOPY to a reserved device
File not found
File creation error
Reading source file(s)...

%1 File(s) copied
F D %1%2
%1\%2
%1
%1%2 (Y/N)?%1\%2 (Y/N)?Invalid switch
0Invalid Path, not all directories/files copied
Overwrite %1%2 (Yes/No/All)?YNAFCopies files (except hidden and system files) and directory trees.

IXCOPY source [destination] [/A | /M] [/D:date] [/P] [/S] [/E] [/V] [/W]
/  source       Specifies the file(s) to copy.
A  destination  Specifies the location and/or name of new files.
=  /A��  �Copies files with the archive attribute set,
./ �  �doesn't change the attribute.
=  /M$ �  �Copies files with the archive attribute set,
1/ �  �turns off the archive attribute.
E  /D:date      Copies files changed on or after the specified date.
C  /Pm �  �Prompts you before creating each destination file.
I  /S9 �  �Copies directories and subdirectories except empty ones.
:  /E? �  �Copies any subdirectories, even if empty.
(  /V0 �  �Verifies each new file.
;  /W �  �Prompts you to press a key before copying.
I  /Y1 �  �Suppresses prompting to confirm you want to overwrite an
+; �  �existing destination file.
E  /-Y" � 
 �Causes prompting to confirm you want to overwrite an
-7 �  �existing destination file.

BThe switch /Y may be preset in the COPYCMD environment variable.
5This may be overridden with /-Y on the command line
�>\������ Extended Error %1�>U�� ��� Parse Error %1�>y���      P�  �þ� �>�G� �&� ���D�s��X� X�rL�>�  t� ���I� ��/
�t(���/=��u���/���� �t������ ��/� �e��  �ێ��C�6���T�\�D�D��D	�D		�D
 � �� ��� �+.�>�u�`�  �ێ����`���t���/�L�� �!�  ���� �ӀB�B���H�Bu�	���K u� �&B��B��b�Bu=�>��v�>� u����\���Kt� ���5�B��&B����+��부>� t3���Ku�& �>����Kt�W ���B��B�D��+�X9at �a&� t�a�]&� �a�g[ÿ��v�>� u����\�[þ����ks�-	r� �� ��>� u
��O�\�E ��Bu%�It� ��  ��� ��&I��&C��Q���S���g9Ys�� ��  � ����g9Yr.�Ct�@�G�E��Cu�) r��@�,�U s�Hu�@��Bt��� �Ct�C����r"� ���S�C� r� �@��
� ÀC�C�rz�>Y�w!�M��ri�g �ra�Ct�@�
�Q����rI�G ����Ct/�g�9[sܡg@9[|�[+g� ������Zr���D�r�Ns �P�]���g9[s�8rd���Bu^&�   �a&� �]�ag�]&� �g)[9[s�[  ��&� >�F&� ��&� &� :� �v� �� � �Ct�Cu�Cu&�  �&�   �&�  �&�  ��&�	 ��&� ��&� ��&� ��&� &� :� ��� �a&� �O&� �)�]&� ��&� ��&� ��H�XÍ6���  �  ���� l�!r	�@�i��H�aÃ>Q u�>S�w�&C���CáO)S�Q ��?�@�]g��3��!r;�t�C��O��H�	��Bt�&B��N�!�s�>�t�� ���O�!��Bt	���=��o���s�B� ���>� u��  �R �B tƀ&B���Bt	��?�����s�B�&>�Ft>�~.t�B ��&B��B t��&B���Ku�Ku�Ku�Ku�� r���" r���* r�B ��&B���� t���Ë�;� s���ù �6��=�6���T�\�D�D�D �D	 �6'�=�T�\�D�D�D �D	 �6�>� t��! ��" �� ����J
P� ��  ��� �0
X�дe�#�!r= =  t���d���R�Bt�o��մ�!ZÀ>� u
��\�� �Ju�Kt����Bt�=��V�;�!s�H �
��>� u
��\�� ���;�!�RP�>i u�P�3Ƀ������c �g��e�&C��g9[r(�[+g� ��9Qv�C�u9Sv�C��CXZ�Q�]�a���@g]r�U+]v�[��[  Y��I&�W��X&9ate�7�s.�>�u[.���S� tg&�&�8& vG�>��6 &�>� u����\��K&���r��&9au	&�B@�� � ��� � � �>��� ���P&���}�&�&B�&�CuG&�>L t &�>D t&�>F u/�>   tV�>  tO�Y&�D�&�F ��
r�&�F��rJ�rH�>   t�>  u'&������� &�&C��\ &�D &�E ��&9at
� ����a�&�Kt� &�Hu�&�H�u�&�a&�W&�]&�Y&�[�Jt���&��u&���&�Ku&�B@t�	���;�!WZ�:�!�	�&�>� u&�>� t�	� �6=�> ��{	�&�H�t��&9WtR� &�a&�W��� � tK&�&�8& v2�>B�6 &�>E u����\�Q&����&9at� ��K �.�>B�K&��뫀>   t�>  u� ��&9at� �&�JÍ �C� �!�C�����!����>D u
�D\�E �B�;�!s�H ���&�Ku�>��6 &�>� u����\��>J�6 ���2��@ �O�\�2���&�Ku/�����s�Q r� �� ��>�u
��O�\�E �J�J�`�]s� r� �� ��>�u
��O�\�E �PV���hsFF��<Ar<Zw�D<:uXFF��^X�� �6 �>=�&�>� t.&�H@t�6 �>��K�� �6��> � &�  ��F&�>� t�� &�H@t�6 �>=��&&�H@t� ��  ��� �5��&�%
� &�'
�&�>G u&�>L t&�>E u&�Ku�� &�G � l� �  �� ����!r&��� &�C��H���&�>� u&�>� t+�ظ D�!� t� ��  ��� �����&� �l � �)� �!���l G� ��� t�<?uG��I��� � �l F���� W�n��SV_� �a[_;�u'�� t�� ��  ��� �	�t���6���T�\�D�D�D �D	 �6'�=�T�\�D�D�D �D	 �6&�>� u� �� �� ��� �zô@&��&�e� �!r; u�=�z�H���&�� � ��  ��� �K�H��A�ôW��	 � �!Ã>i v�i�>�!ôA�!�.�� �9� �!r� � r9R&� �/�!�� ��!Z� �N�!r��.�����Ӵ�!�sg�+R&� �/�!�� ��!Z� �N�!��Ӵ�!�s:��� �H�u
�
 �H�� ��  ��� �l���PSQR�6&���!�� t��&�H��ZY[X���F�uj�>� uc�>� u\�>� uU� �\ ���)� �!�/�=�\ F�� �6�=�|�\�D �D�D �D	 � �� ��� ����߹� �W+���_�WP� ���OX<�t��I��A< u�_�WV�����&��* sGG�� �tO�\�uW^N������u��&� ��@�^_�V�>m uP� c�!&�6k&�mX&�6k�< t:r:Dw�������^�W3ɬ��
w0��s< u� +�� ��A�< u� ���uP�.�X�A�ʰ �_ô�!&�J�&�Jt�T�;�!&�&J��&�J�t� .�!&�Jt-&�����&��&:t&�Jt��;�!���;�!&�Jt�T�;�!&�Jt���;�!�&�> v&�Ku&�>� u� ú��;�!&���6��G�!���;�!���:�!����&�&�> w��SQR&�� &�&�6&���s ZY[�PSQR&�� &�&�6&���s ZY[X�PSQ��Y�  �!&�� &�Hu"&�Hu"&�Hu"&�HuC&�H u@�~�� � �v�� � �n= u� &�&�  &��&� �j��J�Y �E�T �@P�6���T�\�D�D�D �D	 �  &�&� &��&� �"�X� �����&��  �Y[X��= t+= t+= t+=  t+=! t+= t+= t+=A t=R t&�뽸 �!� �� �� �� �� �� �� &�&�  &��&� ���P��������� ���=�6���T�\�D�D�D �D	 �6'�=�T�\�D�D�D �D	 &�>� u�6'�D�  &� ��6� &� &�&��&� ��X�&�����&�%
&�'
�����P�$ &�&�  &��&� ���X����&�>L u�� C� �!s��ڻ ���  ���E�6�DJ�\�D�D�D �D	 �6'�\�T�D�D�D �D	 �6�% � ��� �=�3۸�!< t�<tG�؊и e�!.:�t.:�t.:�uՊ�S�� ��.���@� � ���!�@.���![묀� t��׸ e�!R� &�&�  &��&� ��Z.:�t.:�t&�L &�G� ����.�>b% u7�.��<t@< t<�  �َ�YYY<t<t	&�� ���.�b%&�� ��  �َ�YYY&�� ��ϯ�  �=  t
� ��F��9�r
�|
��	��6��	��� �>�  t�|��F�u��	��	���������F�t^��#t��t���  ��u� ��(�� �KH�6�T�\�D �D�D �D	 � ������ ������sC��F�u0��F�= u� � �= u� �# �= u���� � �
��F@t�	 �$�>�  u0���F�u�$ �� �?��F�u�7� �>��B��6��>E���K�t)P� ��  ������� �� ��Xú ��F����wHuH.�6K>�|:u�&�PH�>�D���>�D&�>wHu#S3��C��< u��A[r&��F�	� &��F��Q��HuH.�6S>�|:u�&�OH�>5E���>5E&�>Hu#S3��C��< u��� [r&��F�	� &��F������Ft� �>�D�H��6�D�>�� ��Ft� �>5E�-��65E�>J� ���� t��I��Í>��6���Ft�` ����r�< t�<\u�| t�- �>J�6J��Ft�4 ����r�< t�<\u�| t� ð W��_II�ـ9\t�A\�A ����s��r� �� �
��O�\�E �SWV�<\uK��?���^_[��L� &�, �6�F� �Z r�A rG&�$�<Yu�L Î &� ��&; u�3�� �c��u�&�=oxu�&�} u���&�= t&�=/tG������3�2�&�= tQV�^Yt	Q� ��Y�����Á>�H�Hu��F�/�� ��  �� ���H.�>�>t�&�}Su��F�K .�l> �� &�}Au.�`> �Kt�&K��K�� &�}Mu.�f> �Kt�&K��K� &�}Pu.�i> �K�B� &�}Eu��F.�c> �K��F�K �y&�}Vu.�o> �T�!< ud�.�!�J��X&�}Yu.�u> .�x> �L �>&�}-u&�}Yu.�u> .�x> �L��K�.�r> ���4 �K.��> ��,�  ��� �3��>?t�����4 s��F@��F��%.��>-����2�.��>�����2�.��>£� �ô*�!QR�+.��>.�6�>.��>�!ZY
��u��+�!���Fu��Fu
� ��F��p���6W��J��Fu	�6���P��D�;�!r���6��t�9��D������D�;�!r�>� t���6��K��F���� ��F���F�t�c�Jt�T�;�!���6���J��Fu	�6���4�5E�;�!s�H ��F�u ���6����>�F t� �6�F�>�� ���F�u���F�u�Jt���;�!Í65E�: ��F�u
� �5E� ��WV_���<�sGG��� �tO�\�tO�:�t��OW^_���< u	�.F� �H�<\uCF����r9�<\u
� ��F�� �<.uF����r�<.t�<\t� ��F��R���;�!Z��R�����1�Z�< t�<:u� �+ �(� �;�!r�\F���O��ڴ9�!r���
 ��F�ô;�!r�o�5E��F�H�>�F u�[�)�6�F� �l � �!< u7� ��F;�Fu#��F�9�!r��;�!��F ��
 ��F����F���F ����Fø =���!r9�ظ D�!� t(P� ��  � ���G�X�� ��F���>�!�P� �6�F�>�F�2�� ���ӭ�� u� &��F��� u� &��F�6��F�T�\�D�D�D �D	 � �� �����F� ��  � ��!e��F� �!��F;�Ft;�Ft�XË����s����< t	V� ���^�.�D �� ��������< u�\�D ��y �Jtq��E� �q�ѿF�i�;�r]�F��EIJ��� uG�� u�K u�Kt
� ��F���H@�!�K u�Kt�=\t�}�\u� ��F����uIJ��VW����E�`�!��Es��W���F�`�!�Fs��_�'r�J�
 u�J_^ætÀ|� u���� �l F�>�� �àPH< u��,@��@�����B�T�OH< u��,@��8�u�J@��������ô�!���ôG�!�� ��&� -@�Uøp%Z�]��]�W�[=@s#P� ��  � �����X�� ��Y=�s� ��- �M��M����#%���!��5�$�!.��.���%�$�%�!�WV�u�u���^_���F  ��G�&�G�6�G���F��F  �G  ��F  ��G[]��G|<��G>+��G=;�Is���S&�&:s� [��6�FSWU�G��F u>���r7�=t2�nu��F u��"��FAtN��<=u��FC��sɬ�C��N�6�F� �G&��6G�</t1�<"t��FuP&�G2�9�Fs��F��CC�&�� �f��F �^&�G2�@���&�2��tCS&�� [s?CC����F �3&�G2�@���&�2���@�&�2��tCS&��T [s
CC����F ]_[��F��F�6�F��F��F��P&�� u��F�< u� u��F �P���� X��X���UQ&�O2��t�o	�>s� �����.G�Y]�&�~  tE��EÀ�F���rB�&�F�P�G+��FX�6G�< u#�|�:u��F	 �&�? t&� u��F �	� ����
P���� X��W&��>�F&�&�eP�G&�EX<u
&�U&�M�Y<u&�U�O<t�<t�<u&�U�=<u��F@&�E&�]�+&�u&�]P&�Gt��	&�Gt��� X&�Gt�� _���G P&��uPSRW��F	 ����`�_Z[X�,� t��F  ��>�F	u� t��F  ��>�F	u��f�� �t��F  ��>�F	uP� @t��F  �� �>�F	u;� t��F  ���>�F	u#� t��F  ��>�F	u�  t	��F  �g�>�Gu�>�F u��F	 X�PV�
�t<:u�| u� �	��sFF��^X�VR�Њ��r
�t� ��FF��Z^�<�s<arB<zw>$��:SW�>�G��t�>�G8tPQR�e�»��� ����!ZYX�]�ECC,�&�_[�P��F��&�F��<+t	<-u��FF� X�PQRV3�3�S�
�tB� r92�������h r,�ڋ������[ r�����R r���I rՃ� �? rF�[�%�[��Ft
���҃��� &�w&�< u�������F	 �����^ZYXÜ��Fu�Ýp����<0r<9w,0����PSRW&�&�
�u�����F	 ����?�_Z[X�PURV���|r:����Ft<=u&�~ un���Ft<:u
&�~  uZF�Z&:F u
�tPFE�&:F uCF�E&:F u9FE���F@t&�G  t&�~  t"&� t<:u	&�~  u�< u&�~ :t���6G�^Z]X�PQRVSV� ^��G  ��G  ��G  � r��G
�t� re��G
�t� rY��G
�uR��G��t��G
�uB�ȡ�G
�u9���G��u�����G��G
�u�ȡ�G
�u���ds��l[^������[^�������F	 ZYXÍ6�G�<�t�RP� 8���!XZ�QR3Ɋ
�t;�>�G t��u<:t0<.t,�<-t&</t"<.t�A�r� ��
 ���u�r�F뿊���F�����ZY�PQRVSV���D^u�� ��G  ��G  ��G  ��G  ��G��w�rS��G
�tU�k�rG��G
�tI��]�r9��G
�u/��Fu4�6�F�|�,u*�D�.��F  ��F��G�&�G�6�G����"�rX��G
�uQ��G
�uJ��Ft<w?u2���Ft<tr,<w(�С�G
�u��G
�u�ȡ�G
�u��[^������[^�������F	 ��G ZYX�PV�F
�u��D� <pt<at<mu N�D� <pt<at	���F���F�D� ^X�PWV�>�F�
�t�W u ��G^� _�9^� _&� u-��F �%XV�
�t�* t�[sGFGF���F� G�>�F^_X� t	P������X�SQ��G�	 :tC��AY[�PR�
�t5�r*�|:t&� t�| u <ar<zw,`�д�������F	 ZXì�  t�Q u��F t���FAt	N����N���SQ<t-< t)<
t%&�}r3�&�]��&�9 t3�&�	C&:t��<Y[�SQ��F �&�F�< t6<	t2<,t1< u�< u� F:��&�}r3�&�M�t� C&:t��< Y[â�F��Fu��F :���.G;�t</u�P�G��^�r��W�X���
</u��F@��VS�>�F u%PQRWU3��޸ c�!���]_ZYXt%�6�F��F�6�F��F�< t:r:Dw��FF���[^��MH  �&=  u�MH�6KH�����>�  u$��F�t�� ��>QH�6KH3ҋMH��=��u������ 	 �MS DOS Version 6 (C)Copyright 1981-1994 Microsoft Corp Licensed Material - Property of Microsoft All rights reserved u � �� � + �COPYCMD= � � ��� � ( ��    �    []|<>+=;" � � ��G    VH ;dHmH�H�H�H   wHvH  HvH   �       �        �HvH	/A /E /M /P /S /V /W /Y /-Y    �HvH/D     �HvH/? �      �� �  �������������   b   �RB��� �  ��� ��O����P�4 PˌÌ�H�؎�� � ���G����H��� ��������+�s��+�����ڋ������+�s��+�����¬��N���F��$�<�u���<�um�¨t��2� �3ҭ�����Î�������t&��� �t�� �܌�@����&H����Ë> �6
 � - �؎��  ��֋����.�/�@� � �ʎں�!��L�!Packed file is corrupt �H��@0�0V11                              �.�/�@� � �ʎں�!��L�!Packed file is corrupt                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              LN   : nN   qbasic.hlp        F          I3  I7          A� I7  �8  (;  �=  �A  eD  �E  �G   K  N  SP   Q  rR  �S  �X  �\  �_  Ng  pk  �n  �o  ,q  'r  s  �t  �y  {  @�  �  x�  �  S�  W�  �  >�  �  �  �  2�  ё  	�  Ô  ^�  m�  2�  ��  �  ��  ��  K�  ٤  ��  �  R�  ��  �  ��  Z�  (�  O�  ]�  ��  �  ��  }�  ��  ��  ��  �  5�  ��  ��  ��  ��  v�  �  �  B�  ��  ��  g�  W�  ��  ��  ��  �  |�  4�  R�  ��  ] � r � � �
 
 �  m � X  � �  # � � 4  6! �# �% 1) �+ y- �. 1  3 [5 .6 c8 L: �; /= l? �A D RG �H J ]K L �M �O �P �R �T �V rX vY [ �\ |^ ` �a mc _e  g �h �k �l 0n �n �o �p �s ^t `u hv nw �x Tz �{ �| �} �~ � � C� _� � z� N� m� �� �� Ď � P� � "� �� ;� �� m� O� Щ |� �� �� � �� �� �� � �� 3� �� � ˴ a� �� �� r� �� g� � �� � j� �� $� ӽ G� �� !� n� � t� �� �� � �� �� I� � �� 4� �� �� �� �� �� ;� �� �� �� �� �� �� L� � Y� !� �� � y� �� �� 5� �� �� �� V� � �� �� �� &� �� 5� y� �� ]� �� 1� o� �� *� �� F� �� )� k� �� � _� �� �� b� �� 
� >� �� �� �� /� �� 4� �� 9� w� �� � e� J� �� �� w� V� �� |� � �� (� �� *� o� �� � 8� o� �� u� �� @� �� �� Q� �� �� �� s� @� �� �� 
� 8� [� |� � E� �� /� U� |� �� � N� �� ^� �� �� #� V� �� %� X� �� � (� �� 1� h� � F� �� �� 9� �� �� *� R� �� � A� h.pg1 -9995 -9998 -9996 .cccp UsingHelpSyntax qbas.exe .fun.character.set .sk .dk .vk .hk .fk .vd .kbsct .rtect .lqb .lim.nsn beyqb ALIAS EVENT LOCAL BYVAL $INCLUDE SADD SETMEM CDECL Int86 Interrupt SIGNAL COMMAND$ Int86X InterruptX UEVENT AUTO NEW CONT LLIST RENUM LOAD SAVE DELETE MERGE USR EDIT MOTOR BLOAD BSAVE CHDIR MKDIR RMDIR FILES CLOSE EOF ERDEV ERDEV$ FIELD FILEATTR FREEFILE GET PUT INPUT$ IOCTL IOCTL$ LOC LOCK UNLOCK LOF LSET RSET NAME OPEN APPEND BINARY OUTPUT RANDOM ACCESS .openalt RESET SEEK WRITE AS BEEP CLS INKEY$ INP OUT INPUT LIST KEY KILL LOCATE CSRLIN POS LPOS .opcom .penf PLAY PMAP POINT PRESET PSET PRINT LPRINT .zpu .lprintu SOUND SPC STICK TAB .vupri WAIT WIDTH WINDOW USING CIRCLE COLOR DRAW .ggx .pgfx LINE PAINT PALETTE PCOPY SCREEN VIEW ABS SGN ASC CHR$ ATN COS SIN TAN CDBL CSNG CINT CLNG .datef DATE$ EXP LOG FIX INT RANDOMIZE RND SQR .tmf TIME$ MOD CONST DECLARE ANY DEF ENVIRON ENVIRON$ FUNCTION SHELL SUB COM .ketv .kbflags PEN .playf .playev .strigf STRIG .timerf TIMER ON OFF $STATIC $DYNAMIC COMMON DATA READ RESTORE DEFINT DEFLNG DEFSNG DEFDBL DEFSTR DIM REDIM ERASE LBOUND UBOUND LET OPTION BASE REM SHARED STATIC SWAP TYPE INTEGER LONG SINGLE DOUBLE STRING CALL ABSOLUTE CHAIN DO LOOP UNTIL END EXIT FOR GOSUB RETURN GOTO THEN ELSE ELSEIF ENDIF IF .ongo RUN SELECT CASE IS SLEEP STOP SYSTEM TRON TROFF wend WHILE AND EQV IMP NOT OR XOR NEXT STEP TO CLEAR SEG FRE HEX$ OCT$ INSTR LCASE$ UCASE$ LEFT$ RIGHT$ LEN LTRIM$ RTRIM$ MID$ CVI CVS CVL CVD MKL$ MKI$ MKS$ MKD$ MKDMBF$ MKSMBF$ CVDMBF CVSMBF PEEK POKE SPACE$ STR$ VAL STRING$ VARSEG VARPTR VARPTR$ ERL ERR ERROR .onerr RESUME errhand.ex -9997 -916 -917 -902 -904 -912 -911 -908 -907 -909 -913 -367 m.f m.e m.v m.s m.r m.d m.o m.h -288 -289 -291 -292 -297 -299 -302 -303 -305 -304 -306 -307 -308 -310 -312 -315 -318 -317 -320 -321 -322 -327 -328 -334 -336 -337 -339 -340 -341 -343 -345 -346 -347 -348 -351 -9999 -2001 -1 -2002 -2 -2003 -3 -2004 -4 -2005 -5 -2006 -6 -2007 -7 -2008 -8 -2009 -9 -10 -2010 -2011 -11 -2012 -12 -2013 -13 -2014 -14 -2016 -16 -2017 -18 -17 -35 -2077 -77 -2039 -39 -2018 -2019 -19 -2020 -20 -24 -2024 -25 -2025 -26 -2026 -2027 -27 -2029 -29 -2030 -30 -2033 -33 -2035 -2037 -37 -2038 -38 -2040 -40 -2050 -50 -2051 -51 -2052 -52 -53 -2053 -2054 -54 -2055 -55 -2056 -56 -57 -2057 -2058 -58 -2059 -59 -61 -2061 -2062 -62 -2063 -63 -64 -2064 -67 -2067 -68 -2068 -2069 -69 -70 -2070 -71 -2071 -72 -2072 -2073 -73 -2074 -74 -75 -2075 -76 -2076 -128 -209 -213 -215 -216 -217 -218 -219 -222 -245 -246 -254 -255 -256 -264 -265 -270 -271 -272 -273 -131 -132 -133 -134 -135 -136 -137 -163 -164 -165 -166 -167 -169 -170 -171 -172 -173 -174 -175 -176 -179 -180 -181 -182 -183 -184 -185 -186 -187 -188 -189 -190 -191 -192 -193 -194 -195 -196 -197 -198 -200 -201 -202 -203 -204 -206 -207 MSG_ForIndexInUse MSG_TypeTooLarge h.pg$           	 
                                                 ! " # # $ % % & ' ' ( ) ) * + , , , , - . / 0 1 2 3 4 5 6 6 7 8 8 9 : : : ; < = > ? @ A A B B C C E F G H I J K L M N O Q R R T U V W X [ \ \ ] ] ^ ^ ^ ^ _ _ ` ` a a b b c c d d e f f g h i i j k k l m n o p q r s t u v w x y z { { | } } } ~ ~ ~ ~ ~   � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �   		

 !""#$%%&&''()*+,-./00123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmm$DYNAMIC$STATIC10019922002553204Use64064K79769313486231D7The7You8Each940656458412465D9The9UseABSOLUTEACCESSAPPENDASCIIAdaptersAlsoAltAnyArrayArrow
Assignment	Attribute
AttributesBASBASEBASICBASICABINARYBLOADBSAVEBack
BackgroundBasic	BeginningBinaryBooleanBranches
BreakpointBreakpointsCALLCASECHAINCHDIRCHR$CINTCIRCLECLEARCLNGCLOSECLSCOLORCOMCOMMONCONSTCSNGCSRLINCVDMBFCVSMBFCancelCapsChange	Character
CharactersCheckChooseClearsClick	ClipboardCodeCodesColorCommandCompatibilityComputerContentsContinue
ConvertingCorporationCtrlCurrentDATDATADATE$DECLAREDEFDEFtypeDIMDOSDOUBLEDRAWDataDecimalDeclaresDefinedDefinesDelete
DeterminesDeviceDialogDifferencesDisablesDisplayDivisionDoubleDownDrawsDrivesEGAELSEENDENDIFENVIRONENVIRON$EOFERASEERDEVERDEV$ERLERRERROREXITEachEitherEnablesEndsEnterErrorEscEventEventsExampleExecuteExitsFIELDFILEATTRFILESFORFREEFILEFUNCTIONFileFindForFunction	FunctionsGETGOSUBGOTOGraphicsGuideHandlerHelpHerculesHighINKEY$INPUTINPUT$INTEGERIOCTLIOCTL$	ImmediateIndex	IndicatesInsInsertIntegerKEYKILLKeyboardKeysKeywordKeywordsLBOUNDLCASE$LEFT$LENLINELISTLOCLOCATELOCKLONGLOOPLPRINTLPT1LReturnsLSETLTRIM$LeftLightLimitsLineLockLogicalLower	LowercaseMCGAMID$MKDIRMKDMBF$MKSMBF$MakeMaximum	MicrosoftModesMoveMovesMusic$MyClassNAMENEXTNameNextNumberOFFOPENOPTIONOUTPUTOlivettiOneOpenOpensOperator	OperatorsOptionalOutputPAINTPALETTEPEEKPENPLAYPMAPPOINTPOKEPRESETPRINTPSETPUTPastePathPersonalPlaysPositionPressPrintPrints	ProcedureProgrammingProgramsQBASICQBasicRANDOM	RANDOMIZEREADREDIMREMREMLINERESTORERESUMERETURNRIGHT$RMDIRRNDRSETRTRIM$RUNRead	RecBufferReduce	ReferenceRepeatResumesReturnsRightSCREENSEEKSEGSELECTSHAREDSHELLSINGLESLEEPSPACE$STATICSTEPSTICKSTOPSTRIGSTRINGSTRING$SUBSUBsSYSTEMSaveScreenSearchSeeSelect
SequentialSetSetsShiftSingle	Specifies	Statement
StatementsStatus%StepStringSuspendsSwitchSyntaxTESTTHENTIME$TIMERTYPETabTheThenThisTimeToggleTrappingTurnsTypeUBOUNDUCASE$UNLOCKUNTILUSINGUnsupportedUpperUseUsingVARPTRVARPTR$VARSEGVGAVIEWValidValueValuesVariableVersionViewViewportVisualWAITWENDWHILEWIDTHWINDOWWRITEWhenWindowWordWordStarXORYesYouaboutaboveaccessactivateactiveadapteraddressafteragain	agreementall	allocatedallowedallowsalreadyalsoalwaysamountandangleanotheranyappearsareareaargumentargumentlist	arguments
arithmeticarray	arraynamearraysassignassignedassignments
associatedattached	attempted
attempting	attribute
attribute%
attributesautomatically	available
backgroundbackground%becausebeenbeforebegin	beginningbeginsbeingbetterbetweenbinarybitbitsblankblockborderborder%
bottomrow%boundboxbracketsbranches
breakpointbreakpointsbufferbuttonbytebytescallcalledcallingcallscancannotcapturedcausedchangechangedchanges	character
characterscheckcheckingchoosechosecircleclauseclearsclickclosecodecolorcolor%colorscolumncolumn%columns%combinationcommandcommandscommandstring$commascommentcommunicationscompatibility
compatiblecompletecomputer	condition
conditionsconsistconstantconstantname	constantscontain
containingcontainscontentscontinuecontrolconvertconverts
coordinatecoordinatescopycorrect	correctlycorrespondingcountercreatecreatedcurrent	currentlycursordata	debuggingdeclarationdeclarativedeclaredeclareddeclaresdefaultdefinedefined
definitiondegreesdeletedepend	dependingdesireddestinationpage%	determine
determineddevicedialog	different	dimension
dimension%dimensioned
dimensions	directiondirectories	directorydisablesdiskdisplay	displayeddisplaysdoesdoubledowndrawingdrivedriverdynamiceachediteffecteitherelementelementnameelementsenabledenablesenclosedencountered
encountersendenteredentireentriesenvironment
equivalenterrorevent
everythingexampleexceeds
executableexecuteexecuted	executionexisting	expressed
expressionexpression%expression1expression2expressionlistexpressionlist2expressionsextendedfalsefieldfieldwidth%filefile$filenamefilenum%filenumber%files	filespec$fillfindfirstfixed	followingfollowsfor
foregroundforeground%formformatformatstring$	formattedformulafound	frequencyfromfunction	functionsgenerate	generated	generates	generatorgetgraphicshandlinghardwarehashavehelpherehexadecimal	highlighthighlighted
identifier
identifiesillegalillustratesimageimmediatelyinclude	includingincreaseindexindex%indicate	indicated
indicatinginformationinputinsertinsertedinsertsinsideintegerintegers	intensity	interfaceinternalintoitemitemsjoystickkeykeyboardkeyskeywordkeywordslabellanguagelargelargestlastleadingleftlengthlength%letterletterrangeletterslevellightlinelineslistliteralloadlocallocationlogicallonglooplower	lowercasemademakemanymatchmatchedmatchesmatchingmaymeansmemorymenumenusmetacommandsmillisecondsmismatchmissing
misspelledmodemodesmodulemonitor
monochromemoremostmousemovemovementmovesmultiplemusicmustnBadnCannotnChangenDevice
nDuplicatenENDnIdentifiernIllegalnOPENnOut
nProcedurenQBasicnSyntaxnUsingnamenamesnegativenetworknewnextnonzeronotnotenotesnumbernumbersnumericoccuroccurred
occurrenceoccursoctaveoffsetoffset%omitomittedonceoneonlyopenopened	operating	operation
operationsoperator	operatorsoptionoptionaloptionsother	otherwiseoutputoutsideoverflowpagepages	parameterparameterlist
parametersparenthesesparitypartpassedpath	pathname$patternpausepenper	performedperiod	permittedphysicalpixelplaceplaceholderspointpointerportpositionpossibleprecedepreceded	preceding	precisionpresspressedprevious
previouslyprintprinterprints	procedure
procedures	processedprogramprogrammingprogramspromptprovideprovidesqueuelimit%	quotationradiansrandomrangereadreadingreadsreceiverecentreclen%	recognizerecordrecordnumberrecordsrecordvariable1recordvariable2	rectangle	referencereferredrefers
registered
relationalrelativeremainsremarkremoverenamereplacereplacementrepresentationrequiredrequires
resolutionrestartresumereturnreturnedreturnsrightroutinerowrunrunningsamesavesavedscreensearchsearches	searchingsecondsecondssegmentselectselected	sensitive	separated
sequentialsetsetsseveralsharedsincesinglesizesmallersoftwaresomesound
sourcefilespacespacesspecialspecific	specified	specifiesspecifystackstartstart%startcoordinatestartingstarts	statementstatementblock
statementsstaticstatusstepstillstopstoragestoredstringstring$stringexpression$stringexpression1$stringexpression2$stringsstringvariable$	structure
structuressubdirectory
subroutine	subscript
subscripts
subsequent	substringsuchsuffixsuffixessupport	supportedsupportssure	suspendedsuspendssymbolsymbolicsyntaxsystemtableterminatingtestexpressiontextthanthatthethemthentheretheythisthroughtimetimeouttimertootopictopicstoprow%	trademarktrailingtrappingtriggertrueturntwotypeunavailable	unchangeduniqueunitsunlessuntilupperuseuseduserusesusingusuallyvalidvaluevaluesvariable	variable$variablelistvariablename	variablesverifyversionversionsvideoviewviewportwantwaswaywhenwheneverwherewhetherwhichwhilewhitewhosewildcardwillwindowwindowswithwithinwithoutwordwritewriteswrittenyouyourzero���ͼ���ͻ�� � f 4   )�   �ր��7�2 $ ��0 * ��. ��_���d F < [�@ <�D Ҁ��N L 
�R�V T W���Z ��^ ��b ����,�v l s�p f�t m�!�� � � � ��8�� � � � ိ�j�� �Z�Ā�� � � � � � h�� � ��`���T�(�e�� t�� � ��I�� � ��� � �� � ۀ����3�� �� � � �� G�� ���� K�S��NL�J0���V�v�.("��&̀��,ꀲ�Q�4B�<:����DBӀ��H~���i��fT�dZ1�b`���p�a�����zxv����ڀ~}�����ʀ��5�:�n���:4�����/�X��H�P��b���π� ��������A���w�؀�������U���ԀЀ���u�����΀ ����ƀ�����ɀˀ���;�2$=�0*��.�������8���xjLJHE�#�d�\ZXVހ^���'�`C�hf������n�vtL�	�-�|.���"��&���������߀��q��D�6� �|b������x���Y�À���������2��+��̀k����>�����|�ـ�� �����Ȁ���������M�0��<%�O�*(��{�&$���]�.9�2��:8����\�HBc�F�*�`N�R��ZXz�܀^Հ��N�vho�l��tr�$�l�z���������@��р������������g�r������耸�ŀ݀��y�����ǀ���׀��?���4��J�������������F���� �  /����xn��!@MH�3Hc����g/,�Kc��oҷAO��R�U�\���7�����A��RiQ{�q�H����,r��E���h��֕�7ڴ�+�x��K. �xqi�~�c�Q���iHa-ZC+�x���f�?c�iJk����S\]��V�G��.��9�b���7��e����qx)4��"�%���z��ÁW}A�p�
���)4�\W�Rý��I�G� $�p�WQ#F+��?b"VP��+�X4�M?�jÈ	;d&ŷQrQ���
���`���!�e+.r�����iPE@K�O؄�N�\��b7I��Ⲟ�˜�,M&�d�$`޲R0oo��`j��{Cw�+�J��q�V�fyFħ�R@ $퐘�� ��7�̈�YGJ�Ue+)U�&��H�)�'��
}�m�����#Rf�I��X`��H.����i[�E�j�iHa.�JÂ��[�)ֈ2J�f�f���,�Rˈ$�� O��,p
=�x�ҢZT��8. iQB����~��+���0��&i4��~ŃF��G����R�O/�����W��:p*�԰���~��f��c��o�m+{HQ�iR=�g�Ґ�������4���7���PP*)|>O�'��F ,p?�<����_���7�ǀ���77듰����jX`V��Ë�Lg���ҷ2���/׬�8�+I�C#�x���Ҥ{��)���f�84��#���x\.��W�\Q�3I�c���5qn�{h����/���A���H��@@���D���@�8��ZL���X
崭�-K	 �cA�4�u�c��E�q��0+H0-��X�[h�|>O�TKJ��v�R��m�,pi��!��,p^�ZU��m"�%i3I��v*+�=9=��&���ʆ�`;f��FK�#�&���X8/m�+홹�!�Jm&�/U���rQ��'l�2�@I�!0	=&&o	�"V}iU�8��VP�˜'��
}�m�4�0��u�E���\_9>Z ��|>r�"�L %���Bln�i��ߖ;S7�@����� �&�M0D&����s�)�\֘�&�O2,=����L %���D��_�f�lYi��@E�����&|!6	��D&��eeU�Ǭ���!õ�dy;Y�i���E���a6��L %����3�	�e��D&��Ⲑ²�"��E���;Y�i���r\V�����a�L4�z�"�����<	�M�m3"!5�������5�h���q��ޞ�k0��v�L !�τ&�4�4C�eU�5���v� ���"|�e����"�L %Ѓ	��&��G�ǋ� ��ZM��C
˚�1%n�`a]�$�M��0�A(�g	��O�Me!�e!�e!z˚�1�=�&�f����j�����4�L !Y�wk8M��?�!5�)�QeYHaYs[Ѓ�kA #���@K��+u����h�	�Blt�0�����/�#�f��ز��"YH|��=e Ee�i�!����!õ��@K���Л�a�r\�վ���"��2<;��q��D&��²�Ⲑee�l�7k
(��f��B:&	�W��� �M��B�5��A���i���j\K�"Bl#ND&��*˚�p�c����!H�R ��Ɖr\�վ���"��2<;�2�@I�!0	=&&o	�*������VR�(Mȇ�S�N#��>�-P��!�&i`Qph,. � k�Y��N�jv�>����\M��/[���S�ƀ
��Pv��� ���f�;E�4�q����*(�i 5���X����fc�}�x,��/f�ӴZ��n���������ÂJE��������EĽgfe�F!�P��^�>�厤ƀ
�<���Ke�Y��
��$33,r����W]�t��
�?@>�Q�xg�NÀX�(�(�x�/�4�^�_ϲ��� ���n�������)�)m��Ǘ݀v҃�^x3�xH� �t�w�f��D:���8F�s����lg����;���9
<�@5қ��,H�!灀�dC� ��+�m����f��
)�r��_�:���o��J���;�������!�{��f�Կ���i.w��!��ƿw��>�A�^uqiv�EӴZ�o���z�����u�z�\]�}i������u������Ո�Ǫ���,~��V�4���?�r\�վ���x�<ߋpV��ůe��`;n�n�yZL� &?|�'�t�X��������}5��T��o�i3H2�?W�3x��-d�����J��S��SK�u�pjX>���T鈱5�H2�_�J��zD?]����B�"���	CH2��M��v�Z7��,�"��n��p�5,u��I���鈻RA���K�×+I�C ��.�Y�H�i����ve�M�6�ߊ1��{b�����߂侙A����\�.K锑H����&��}Ar_L��@~OyZL� >;;	�M5����C�{c=�E�<�I�Lh���,�$�4���+���Ml.)
��"۾��!��ȶ��=�i3I ������[/�iD<T*��UZL�,�.xY�H�i�����-�8�ҋ]�E&��=�i ����k��m�t�P	;d&'��� $��3"%VQҲ�YC��Ue	���6Jw	��u;�E�|�0�0	��L�ԣ����t�DrJY�����.����T&>�,�ˮ�q�_PiVʰ��'��C��/�D[ui3H� ����t�D��̀��%"���W_��IB��Y4�e[����IH`�q���R��]F���כXk���R,��_̓t�u�v	����Z��61�Q!������7N�#��+�m�c�0�-x�H�0W�X�����J�f�r���Lt��n��SB�H<]v���������Y��3ߗa���큞���=�XM����/� [���r샀_�@3ߗa��'��Y��:�� ����P�B����e���*G�ҭ�5�iW����]v�"���v�.�	mդ� �G����*��t{�c�12��B��~;m���6((�S�;MWX_P��"��j��M�G݁�͑���ԋ�3�d�n���ZL��F�-6-{võ��B��~;m���6((�S�;;�:��vf:�ݩ-AV��Q�����w8��Z�&(*�p��Z����6�}���RV
�f���o���E��TK~�$&����xZt����Ď�D��_�f�@ $퐘�� ��7�̈�YGJ�Ue+)U�&��H�)�'��
}�m�H/�Ң��dj+�r�_PiV��X7����A�V�4� :m�Hg����_�f��8:�UU��N�w� ph����@�x��~?O��� �H~�b�-J�u�)�[	"�!���Y�V�����5ՁI����q��5ՁJ�e`���F�w�nS�T��XKJ���|E`V���E:�IVL_�W�֥���!���~ʰ�4�V��r�ZE�Ң�1_4�1Y�ƞ݃J�� ��WqJ��+I�C�{���a$i5��x�*ŤZS]���&(oY)4�F�	5�}/]K���J��W�`2)l[q󬝞
�۝qc���%�����"J������
bRZ�}�2�@I�!0	=&&o	�*������VR�(Mȇ�S�N#��>�-P��!� �Ay�D>v�\.4�6�j�f�`Ys�!��	���~Z���{�ٮ�$UV��O���	�x��ƅ��G��	"Ѵ��ZҞ���-+�Z��V�Hpk�`٥Z>�|<��)0������J�>�s0[��أi;�7)�m���$C�!I��u������1�DG�J���x�ʲW5�+�4����kH2��� �D!�U�r���"J�E&+48�~]M)L�I�A���pkJ��4�W�ZU��Z=K	"Mk�����7ڴ��Ɔ���@��|pF�J�o>
�e|K�u,r�+H���}z��״�,V�x!��f���Ri\II�}�r���Ɓ� Oهi4��aIV|K�u,r�+I���<��԰iQ?jC�4/����uդ������0��R@ $퐘�� ��7�̈�YGJ�Ue+)U�&��H�)�'��
}�m�H7��w�
�w�`��^��!w_���iQ��~ѩ3H�9���MA��_��oz�A��ƚ����5���j05������jw��3P`bf���ͮi �5����Q۳1�JkaqR����~&�E�?�X#�AAo_`ҭ��	 ̾�B��]�wy���c�Y����������@SZ�t�*Oko,�\�@���"������GKx���}(�Şv*t�X!w/׬Ա�����c�̑�ԛ�D�����Y&�/���~��&i1A��`�=�jX<J/I�� .q�`�9;�w�I�a���#s�X�ðI�c��d[v1�5�8������0\)4�G{l�[���װ�Qa���"qJ�g�7�JE�x�^�]������J/���C����pkJ��Pj�(;n�	 ̣i"�-�C�to�ү�hpkJ�f�e���L��i^��t�t��}@_B�T���Hea+I�E�?Ζ��25��V�f\MqQW�.m�Oso(�L\B���6t�Q)KGm&���_��4��;	�Չ�X�)0�M}ZL�b���������AAo_`ҭ��	 ^F�S�iݿ�y���az*��z���֌k��e$R Q$��� �Gڴ���M�)����E�԰��7���X
|RRb��qo�4c��kc�}J��+��� ��5�W�o��@8�h�Ҿ=���&i����a+��wMKO��m]�UE�H�a|�!�Y�������!tB����v�LOG	�@I��fDJ���e*�����Ys$l����w�>�T6��aH`Q ~����i|�a!D��Gݵ��/ɹ�c��$X1?�R \f���V!����8$X���R�� �t��lz'"��_N�~Abl{Ӵ�Y� ��5&i1X�|��9/���׭�ݻ��AI��0�k/�!���Ӥ�c���q,`�`�P�q8�2zt��p� ) 	���1X฾r/��&+#I0)5��B���|�8� ��G�$��vHQ��h)1X� d :<kd�E�rkaq��t�4�@��zv�P���T��z��4�1X� � t�'�û�0M00 丵YG`G:�s��N�&+4��t����N���N��%m�aL���b��L��آMl.)
 U���8� � �r\Z�,��#���l'N��l��������c���%m�aL���b��L � Ǝ�Mv[F��4�# bm) �5۰�{�MvXc��&+4� �û�3�06J�v�^���@n��'N��`
���=��00� G��VطN��`����[Fq��� �2��Ȟ$������ٙc�Ӥ�c��� #���Y݅�[����^��w��v�����-:LV8i�W��C3ò�;��`�LM����F6�i�b��Lw /ϲ�qkd��\A��b�06J����.�^5^�:LV8i�W��P$�Qc��A�k��t�4�+o�}����t�1X฾r� \_9:� �#E��,v�o��㧦A�ZC(�� ����`f��(�YJ���e*���\�%;��B:���O���rR #��D<���� G�;m��>rB�R 4�k����hH���.^5���z��O�i� 4��,r�l	�y��y"``�x�5,��8;��o9����:C���Ȧv�4�r�4��}b�4*;�!�>���!��O��L��`i���Z���Ht ��u,8:�����Q� b`��"�ڤ: i�x$����v�o9��4�#��r�["|���
C��7����俉x�A�� ���c+1��H1:C���X�@�A�i�./��gj�� ��r)���Ggׁ��ȇ�9>Z
C�}=�dCϜ��@����َ0��!�L.�+���)��g� � �=X}FF��Ht ���#0h����X	i1�0�:C���Ȧv�4���-�CHi� #�n��dC����[@��>,�a�t�@06�.���@�0�``@��|XcK9:C��D���C	a� ��r)��E���Ȧv� ���E�x�/������&|)�v�LOG	�@I��fDJ���e*�����Ys$l����w�>�T6��aH4YjTW��}l1��yGR@�SU�+����0��4��U԰�������a��!��C
CH��Z�eRvu�|X�a�I.3�||GHgdC��qo/O"}Vz��i��!Ґ��X�3(�A� 	mSi x�cE���L�R@ $퐘�� ��7�̈�YGJ�Ue+)U�&��H�)�'��
}�m�D/�iV�L��ҷ���c�t��9)@�� Q�/�p|[/�a�>iP ��E|�X�@�0=��
U�\,S��y�|�0�Q6���4����2
A�|�U�V�ƕ�x�
&��`�Hm�e�o�E������x((Xi����1�o9�a,�e(��m'{^��X�9���(x�v3���x/�_�c����Ȟ;�6��aH` \A_��X�]M�<����0ФB���Y.o9���e�
���_��7��y�x�H@Ǎ�υ!�N�	�@I��0	3xLȉU�t��VPⲕYBk.d����p!N���j��9)1B�P�`W�J��mZV����Afrk��%c	a���{m��!�#7�S�d���>٨O�a��jCo�����Ծ����<�%��ACJ��q�aJm<�i�rR�E����`+�#���3�"�D�w��,�#���1�hD\�(������������ȇ�!�c��ʐe-�-K�[h1�k�x&&��C�I���R��6�n��;iM��%R���0���a��yKŎ-�����+홹���Co�����Ң�V�"�#�����yK�~���J�J�Ad@Ҥ{b�A43y�#	t�y1Ɖ~�f�D<	�
C(�� ����`f��(�YJ���e*���\�%;��B:���O���rRf�/�,r��N�j>)��x-D�t��ⳤ�x�S ��J��q)4��=��v�[7��I���]M�<�kd@&�^�4����R��<ݤBo9�aI��ģ?��81e7����+D82W7����P����,�{h��[�qB����sO��v��7�.>x;��o9���%&����+���d&�fu�+��yi1A��8;�n��y�ټ�g�4���\��05���<�<_�b��z�_H�05��7��l��H3-����XϠ�B�0iDf;i;��_P�x�q6�_��9Gc1�I��ׂ�����3���t�'��3I��uX�3YAE�g��A�a��Α�|<Vt�@@�<J3��s��(�	��y��4��������s�� ��y�)4�� �`x�g����c�o9��I���V.������y\�9 �[c��3�o9��<y�)�v�1�ky�/��T�м���<:dxv�d>�������7����ƅ'�1����K},�æAǇl�M�<�<9XФ�'0ol}�`G���>��Q3� �x��-@�4C��<�ks�"�Q�ݝhn���]	�y��y ��
G�_��݊Q43y�7l�Ij[��)	�y ��IF)D�<��8R{B�<J1t&���<y�)=�82��M��x�#�o���b��&��o9��_Nԃ�o���b�LM��s��%�L�b���k���3�������L�H�>+:M ����S�����Q��ų1f�m�H��.Pj<>�XLe`�y�31
G է�G���<,�5,&2��Mʎ���G[��N���<,�5,&2�����I�u԰�_P�����CR�c+0��y�x|��@�ҷ�K�+1��!431
G o����s���`ҷ��2����:� E��.b�הi[�XXC������y0�{-�c�9ټ��y�<>4���:��0�D`�C�j&s�`�&��Q���R�]_PiQ-&-�����y�/�M #��ϔ��J�i0z��C�y�8�M #�J�۽@��ҭ-+{J����y���M #�O��v(`�o9�H�:��M;b����вV&��E� ��cD@��5kzN�
C(�� ����`f��(�YJ���e*���\�%;��B:���O���rRf�~ֲvx2����Y5��h�����~+�G�.K�QŔU�P[��M�UY����'��zUUY�^R?X��*��UV}�RJ���/),R���cUVjK�60UUfu~R�Rߟ7��!K��I�E�(�fQu�A��/���b��|	��	��	�||�_)1�R���O�!ǀ$�����ߞR(1J%���F�Z�f�e������<a���'�x��	�> �?)إ��S����I�Lh��׿�q>og�1��4����)lR�?7O���!�?�����"͊U��������B?<���I�Sg�{�~bx�xs�~x��ϔ��)nɘ��ݯ�s�>w���R���	�&i1@����%7����c������!�����M�� ��,���<g�~.M������x�~R(�K8��&k<-����R/إ�P�>~ �i3H0p����S��O�x��cG�6��"�4x5��)�O���������T��)Hq{�4t����	�~�S�G��:���4?�fl0�&7yH�b��}��GI�m���ɘ�R(�K�(xx)3H���H<�8|��xR�����&>��:�H��x(�]���>�|���R�4�17�^��	����,�K����&u<�f/�7+�Y�J"��l��)xz�^ ��M&)D{�R�]x<y�gI�E�?6/�L����g!@�Pf�Q&�l%���{�\�{��F�g�OC�����6���Y��	�c���?<#�fm��eb�J���11�&����l�x�fRG1Kq�f-&i1B��$�`+����|Gvų��/�J+�{����&v�	Ǿ���R�?7hBi��q�c ���I�Sc ����nS�60	�? ��7�f�)����M�x=��_��:1J#��"�������_)��؊�i
�����-He ���B`z8LL�2"Ue+)U�8��VP�˙#d�p�GS�|)�Z���C
L�cX�>��7�X�0��I�	�x�RC Y���A��0�M^m�&i4�p@�p7�S�l�,���JEZ�fx��� �Ϸ��c0-�	�H�Ç����^x!@	o�����?�I�lN�E	�9`W��v�َ`[��E����ϡ�lN�E(� ����A��1���'M"����V���p`[��E�K���`SA��e�`�t�(��r\]�$Z��T��'M"�v^X��Ű�� �4�,8���|�`[��E�>7�+����lN�Ez�3x݅��T��'M"��;��vd��0;���,��t���y�rJHgf�V5�'-@��4�`Q���x<�!�&iXqq��ϡ�lN�E20@��'M"�7�Hg�I�2kaq3�lN�EMa�C� �4�,8_�Y�_�KjƘ���"���kdC�L�(��f!��j�:�`[��E�
6H<�������۾�m�f�A:iXq3�H�K. �;�p`[��E�G��l�(�0��a�lN�Eh���g<��'M"��D�[c `[��E��c���A� �˘��~���R�$���[����H9�#�k��Qafo;E�
u4}�dC�z�`�t�(��E�������lN�E����`�p1��0x((��#�]Y��`!�����L��c�'�DyVR��5���3�B�	��m
�#DA(�gHe ���B`z8LL�2"Ue+)U�8��VP�˙#d�p�GS�|)�Z���C
C���l<x(�pB� �Cuϐ��`r,����HO+@���8n���e�&��6�����Q�#>`9c�ʀ��8���&� �Lp�,�%)�'2�!������s/�  n^3���:��NFf�����{c��4��1����1�\� R�@��Р�ާ��p9���7/��c�΀��I�q����A@-X�s�z�8�y�����u!� ��@vڟ���Y�!�n^3�����_0���a����\���@1�ri4��%ˎ��'#0$7l^���rzr 7/�����A@
L$�8�lp9P�8��y�R�%�Pi�'1�p��Hc��찅�tR��s���$�;@#��r�i�y���c���a�%���C��ʀ-����rzz7v5��t9�J�Nc�`���Ð1��@-�8K9=�p�/�-ԇ@������݊?����@ �ݶ����s�i�	9���8�Kky��c��� 1�\�H=t�@��`tϽ�a''�0�p�'�8��Cs	9�Pf8����<���c����o��,����@��K7k#��8��>��������Nc� ���� �c��1��%���p�{,��@�g,p�Q��	9=Pc�����#3�20���`������p94��(�	g*�1�Y���!� �\��v��I���s�vݙ�c���@,$�8�F8�G+M2�ݎ� �c��� 5ԇ@�g������NOy���������a�	9P9kf��I�8K9��8K=�ۤ: ��c��1��I��>��y��r3��r�,lp9���M: jc���Ht��Y�pG��@�c0�����Nt@��w�����Vr�z{9���&��.�8K�r1�Y�ZC�̸�1�����Nt%�*�;��NF��a'* 4�s�if8�c��1�\�`[%���I�A��5��^�/.w��7\����y�`&q�j!�'#+	�{���,g�K%�s��_���8K�P�$�X�{,f�Oy��c����e ��e��C��c0�Lp�i��	�˘�/��>�Ne����q�4lp==4��1��g���ea2�A�1�X�88KP9�c����c%�s��ӓЏ8�P��� 4�p=��c�XL�	`k��,f��%�K���#��1�_1�4SNt���{/��t%���ќp):A����=��	c?��lp��z(�	�m��,�r��ӑ�[ke�|����p=��H2��z�,p�3�M��4ʘ�/���8K4�@�Ә�<X�{,�&�� �X�z3��H2��z0]��,fi��`w1�_�0[F8K4���c��ʀ:�p==9c���-�F|��T�+	����	q�!��-B8=%�CM��: u�zs��Oe�����r�p=�BҤXL� �1�\t�qlp���D�	|� U��#05�8���1����{t i���8�1�A��������AI1�Z��h��/�X�%�c��1�������� �lp=���c��t�\)V/C�=8K���c��`>&8K�=S%�T����C�c����U������{z"�ea2�!m�p�3��	j�18K����	f���8˖��������{�i�c��v�� ��e��C|c����R&8K�9~�	|�0468K4��c���y�8���c����#����0?�~��c9`>,p��!��%��1�_4p>p�i4�ұ��^��O oX�z3��8L�0�c3Џ�p���&i �	��� �1.�MgHe ���B`z8LL�2"Ue+)U�8��VP�˙#d�p�GS�|)�Z���C
A���Y+�+	�0�a�=s�a?�b�5g�x��C��Sט���A��d?T��Mvd�[%�=�@�L8"�n���sR?Xq��	l$����1��-�L8K`�8�H�a������_�
,��=b���(�?Xp���	�W�a����[�a��A�e	t�����3a1̕��q�f>�͋L8�6P=�~����%A�����Ўb���(hR?Xp������+�0�ef>����p0P`�@gH�a�'����1Y���ſ�?6P��~����fid��Å�1�9���Á�3�
��n����9b��#c���^���L8X6P��~���8XL�l[�a8L���X��Á���z�9�4�q� ����e��o��钱��-�0�a.[=r�4)4�py�����b��5�4�3=b���Y뗠3�~�����Q�e�ط�Ã��@�X�A�L80x雬b�M#��.Y+�ſ�r���ط�ÌC1Ŕ�?i�8�1e-A�L83gſ�?K���'�]#���R���Å�1�j[�a��(�f-�=�~��~Ŕ�f-�0��f8��L8~y@,pXO�#���,��X��ËVc�����Ìh����_�Α�Í�,�NX��Ãc��,[�a��X�����G��G�ط�Ã�1�X��Å��k��,pG ~(R?Xp�dzzſ�{@���%q�ط�Ë�������G�4��=�b���,p*�\q���q� �,��sR?Xplő�͋L8 X��W�ſ�/�^��~i�8~1d{ſ�]�����pAe���sH�a����	=Pb����C0,p #����Ç��F ,ph0�it��G�X�50���-�0�mg�9A�L8 �,8�=�~��g]���[�a�$��{>�9�ߌ[�a� X�U���6M�b��K��� 6�cE�x�b��=k:C(�� ����`f��(�YJ���e*���\�%;��B:���O���rR~�XI�n��y�� O��6��z�3�A�1�XR�RcB[%d=M����m� ��bױ�ǎ���`̷��n��Y+�����@�ZG�^�)�A�����MI2W� ��m�XbR�3d���P/�M����#�X���i��d�H��a� )���ſ��l[���B��:�
��[�Ԡ���~�#�X��E�Q�����Hw��%f��}C�����v��h��q��a��Z�G݊ W��z�@�6-��x���R=����G����Y)���0�a��:9�H4o��RY���JXg&��W� �Pb�7�ʄ�	rش��Ѩ`kL~�#�������8��\���-�((�y!@Y/X;c=C��Ï�w3�h�=��gz�H�����:����K�ȼ��)!,fŦ��}A������	lZ�gg�ux((��-�a~�]l̾�B���� P=b�(�5	I;���8Ť{	�Z��!^�-�1�@
[k"�4�b�q��f- ��������͋md^qx��ib��GFq� P�b���m��KP=9bۺ7��9����3���<i�z3b�7�8�y~�,Z�/���+����X�\	�{��-#�G��Xc� ~�k�a�6w݅��Ef�ԇx�1iK})�L~�?%�j��� +�;i�����1i�Ơ_P��c� ~�j���;/Y qH��K�y���lY~�?4�a����0�E�h�m����ŗ��fž���3_}��`Z��(Qa���G�c��?#��jM�A�u!�u!��[����Ez8pa���A�HRb�o�@�)�>_�n�qqt��>JC(�� ����`f��(�YJ���e*���\�%;��B:���O���rR/���3�����iR�:lװ�Ң�½6D*"RC�ԙ�7c������_��$'	�8VS����/�;�p��|�$'	�8VS��q	�.�c� d_�F|��&��YH|���}��'�.��a0�a�q/ �	�h�*�<�.f>zA���S��׀$o�dh��)�v�LOG	�@I��fDJ���e*�����Ys$l����w�>�T6��aHw��7�gK"��㦐��O���p�x��r����399�*E�n=��|�P�9�99)�v�4|�P�f�~(sR/�f\C���a���c?�|�(���{䱟�>m|Ԝ�f���~5"���f�[�g
��Oy�t�fOU�9=�4�/�qԊ,p0�y&�[�`������8�<�4����/�:Ԝ�K_p7�R1��_vke�fq-Y��:<�8�1�Ɓ�ΐ����ke�f�3VcՍћ%�?Y�@皐�1ƈ���2�@I�!0	=&&o	�*������VR�(Mȇ�S�N#��>�-P��!�"��Y��&t�+:^:i�R�<pa?]!L�׍����jE8bk&����v�p^<���%���CKF�I�a�
j�GhG��鬿� #D���!�b�@嗗H4FΝ�����.k��a���f.�D��c���=��C�X�=��C��4��8�т�=2l�x��_��|o�ӵga�{��ⴀ$)��_�F|��P	;d&'��� $��3"%VQҲ�YC��Ue	���6Jw	��u;�E�|�0��f�L�dVt�t�.Y��<Ha?�!�<2sY2�4��#D���py0��
sHi$��ǔ�yt��"AqZ?�12V{䱟�>m�K�;���h���Z�����Hi$�M��%�>�l�\�Ni B��w��g��'#=r�C�Hi=�n��y�p7ز��/.���F��B:&He ���B`z8LL�2"Ue+)U�8��VP�˙#d�p�GS�|)�Z���C
LPV�;t��8T[{`Ѿ Ӳ!��ӝK5&i��s�J���l�#�@�]/��?Zs��'�uٯ�D�]v.���0 ?�4���j0��F��ȇ�"*Q�-F )�py�9a7MK�o��#����i3H2���o��`B�P��*�U��H�=Ku���V�4�(�A"����\^Wc�]kR���E��e԰i��Qlg�}�8jԏ�F���*Ӗ�]�vD<T.���zl�,� � S�Q���t�n�!�4d��Y�(8�v� `����#�j5V�4�auf+	��r¾Ϣa0�ɏ����YH6���RV\�f�;�h$>;_1�.���Bp�#ʲ�²�c�C��	��Ek�Ը��D�2�@I�!0	=&&o	�*������VR�(Mȇ�S�N#��>�-P��!�"�.�vDI��cR�?E��f;i5�!����ZLP����N����}첇�l..�Π��-�^K�`��Ը��DV�4��K�5p�m��{�#�Hl{>+������W�=wĐ]��)aFÃs~�;	��E�:/!�_�LE����a��"�MvE ��.��>1I��탦C=��l:��f�e�����i�l��@!t���b��:v�PC:E��H<X;`.ݰ���s��4h��m&�D<T�*�f�e��z��c�ƻFF,8�!����t�X!w:���5�.��锰�a��au'ޢ}�HQ��H2��IIB������}hȺ�)l��j�`�gz����]��!�"}�3�b�:l�Mv�V-�^_�MK݂Pv����f��7�	��S���԰�d0��?o!�_�LE����H`JJXg&�8.��b�^�׋
5X� �Zw_�[(�5,8.�e��A���GŶ*�F�RrDk����GŶ+I�C�.K�Y���LA�Z��l8,�\�B��_%˚����Z�����]A��]kR��iD�˖��F9���:�qv�Q�4����I�������},�ð���I�E8����(��x"�>�@�a��M��!E��ݗ_�FKu����:F��t�I�_�i-X�~
b$`~,x:N���.�cņg�	��>�Cu���'Or�f�L���cX�~
wQ��]�8��E�at�����j��k���&�xj+H�a��f�L����p?5�KP!��Q�/!�_�LE���0}���PQd� 2�í�v���ZA���@�!H�,/!�_�LE�t�iLF���]�5ZH]�^���� �7��,��~
o͵�p;R�]v)���!t+�鈰B)���15�ݵ$f-~�Pb{����mv�Ը�r_L�ƶD<h��%t�?�H�c��)�
�!��Q�/!�_�LE���0}��~�fx�Ƨ��{���ZA���y]
�:b,��F�3�LF����P�3/]Ct�?�H�c��)�BB����.阅���͞5SѨ(�n�x4�C=�[X���Ÿ�ArX�((�p��&5��y]
�:b,��x�˷l;e�0}���q!�z��m�HP��V�4�R�cE{d��C(�� ����`f��(�YJ���e*���\�%;��B:���O���rR�um�cņg��L[�½�6D$jL����g����Z��_�o2W3C{Y�e���:/Δ��8�>v��͒�����f��N#ڊ�=x�X���!�*+��͒�(��Pd�J-v9�SV<��y~a�I���t{0Q)0�(��P1n�Z�8sĦ��L�/��"���Mb`�#�S밯C}� ��4��p���1�~����C��Ս_�e�_�<�JC�.M�7��8��C��񷩋,G�yH�a��>'��9ǖJ����>'����E~�_�/صfl��I�Lh]Y��`!�tL�a0�XW��BDG�e!
�YH6��cܐk���!k�<�%�t�hNDyVRV\�}cv$�#DG,+��)�v�LOG	�@I��fDJ���e*�����Ys$l����w�>�T6��aH���o
b��,\��dAtm�� �DjL�i�^��8�
S�i�Ҧrw�z���1̤�9�Qg�����د���<��դ�&(��a/}��K�@�qm9�+qg���+���%������h���}�mn����W�����I��h�m٘�%5,wau�f�<�B�#0�y��ZA�����W���<߅�E��i�/�Բ��޽���kH��T���.������.�/�4�M�� �9f=�R��@�Rްj�`߹ S�Q��j&rq�g��R��CN�{Y����Ս_�������7g��O�ZL�?BnO �P.���z�������XI))����g&>fqu�C��dr�z*�f�&h���t
���������B���0r֢g2��8�+�Ѩtx�K������A�6Ң�.���[��TQ�k��A��P"�����"͜5�/�4�c�!���5�_E�jXa�"�5}d@Ң��t]��:A�N�k�4��,�~�F��H�`�� s��7�m"����O��T�lfr A՞��f�egQ ��H�Y#�Fˮ��]�S��s�{u��ng�"	U��&�L����A@^?Y�u�U;�t	��D�\1Y��R���n���mN�@j��"�P҈O)Y����?K 6����+I�LP���&4�+#}_쁦�FȀ���~�w�9j&s�Ƴ���f���;��qb��RcY�Ik�u�e��"*�i[���:C�8o) 4�o���Ҷ�Y#�Fˮ�G�ԙ����A�n�� �e�B��֑��><0���+H�go�7�J��M������`y�ی�W����������0�)�������50<����'�L�iϬ�~��z�����_dqu,$:0WŨ�˂�8��q��o(�Y&�Ң���*)��ZA��iD'�3����Q�������G�8i�RN���_PiQM����i��[y��x��� �G���
<�*Ep���ơ)'z������`,wN�� �`� #Rf���c�.�`m�>�9�I���9D}n@{)RX,��Γ4�@���{��?.�ų��^":1��Z���,��c�Կ�_�� ]&���k%�J��0z�l���R��$�5	 ���P҈O�^4�?�W}�a�4�K�

�&i!uf+	��b�3�M��ɏ����YHB�����3�]�����|ǔ��-	�h�*�C
˙��n�c�#E2��B�O�C(�� ����`f��(�YJ���e*���\�%;��B:���O���rRF �f\��v+|d��$AsB/�
�jXHb�I,����H���}�!GǇ�ZL�)�R���q��D!j�6{Q-��q�S0��E�	?-�$�Ne/@R��NH��_P��"�E�Y/ـ����u
�p}�ve�Y��E�5���,�@��X�.-�'ѨHR̤�#�����ŤZs)x*(��W_dC���}C�Q�V�f4"����ܫ�@�Nk��E��G3���m��dC��Е�~�����R�m�E���:��¾��J�GhGUj"���H�a'�u}�����5�����l�vc�9��j*(�_�EV����0�+I�Lm՘�&�$!6y�=8M��B9a_g�	�1�)+��5��P��A��1�A�w�܇���~�����)��'m� �o ��'�!�N�	�@I��0	3xLȉU�t��VPⲕYBk.d����p!N���j��9)4��s[�8�`.xP"�DR}����+I�t�(�z��@�H�#����2_PiQ�!HQK~V�4���1��1�d[n2S&8N�ld�Lp����Ű�Jff�ea'၍��E����J�����R-KZ��+%`"��R-K�Y������^ÌQF��G���"���(_�݄x-D[����	��P��\��u�7�@���N?R��^}Ƣ�,�V��U��"�gdjH|a$[j��1��_���C�N�0�%��c�����I�a3�Ԑ��l�!ާH���#�E
C(�� ����`f��(�YJ���e*���\�%;��B:���O���rR%��`(�X���
�,pp��ZL�H���_�6���|j��Ԫ���L�3H�a'���	���}BH�_H\R�%V�-��4�l$��h�aDCǰ��_HW���yv�&iS;#R:0��Rt0�>�2��сO���I�a$�����#{���C�	#����)�ag`��K��U:O[	��!M��7DR�>��@_K���$��}/���I��H�)�b��܁!J���g�I�IwVb��	=a6&7Bl&z�����M��A
P��&=e+(Me	��5�8��5�&��=��|]���]���ߏ�qn��1ƈ���ZC(�� ����`f��(�YJ���e*���\�%;��B:���O���rR7��^�W�J��/�Hb�[�5�n�o��A�E��$1i!��7>1�/�^V�4�g��%3	�[	?�M�E��D�\b��nF٤YL�H��g�Hn�H��;՟��=$)� /��B�$���pq���6	g4��t��}/����= Xo�G�,7��a$=V�<�I��t�&@ܦ!ެ�50!�#�{���I[	Q6���C���}/���I�G:B�$�Hq.m�g������!�՘�&O�a0f�	���6Bl&Ln��1�(qYBk(�YBk(�YBk(Me�{��9�v�RM��*���T�#D��(��� �]8�He ���B`z8LL�2"Ue+)U�8��VP�˙#d�p�GS�|)�Z���C
LRM��� ��u�}iQ^`�&��@3f��QI��9P �7�iQF���J��n��ZW��i3H�f&Jd�W3\Jeni4�I�]D���.�/�4�^��7Ѩbw�*B��:��Du����o��K��>Ei3I뀓;!1�VRWYs�D'y�7����IǾ��&�`!��N��DLz�:VP��:V\ǰ���k��v���#|B��'l�� $�p���&dD��:VR�(qYJ��5�2F�N�8��p�S�Co���{�AAfrk�`�\+���Ȃ@��b�@\Q
�I�H�7�u�o Q��0RD�Fq�G����x���5���d�4��$�86c��E��D�\b��nF��	?V:]DQ���~K"��IU��r6�a'႒a/`���b�4��W�o�D[��>�&0�&i1XI�z�3,r�5w��i�s�����O������´��YL�I-��7)�4�k��j��S�������q�1�!����/�� ���/8�� G��&i.��a0n/�����L���yBl&	k	��G,+��!?�Lz�:VP��z�(Me	��5��k.c�]��f��ߏ�4'j4����� |fb�@ $퐘�� ��7�̈�YGJ�Ue+)U�&��H�)�'��
}�m�u��\�"}.1U��'D��w������Ka'���	���}BH�_K�UV�-���O�GË�4�\�����R��&�j"���V^�.��_�@�����q�H�˴�����C���4�l���p:��!I��x�1��ⶑ|��d�J)G�i
L��%s�
L�͒�P�e���~fJ��0�z�����l��f�I����.���� |[�4���ZO�/��ei3H����݄�7)�w�?MLzHS{���H|a$s�>;����z�L�)3I.��a0ct'	�c�P�˘�!��~��"�LŤ2�@I�!0	=&&o	�*������VR�(Mȇ�S�N#��>�-P��!�!�⴨���F�}�qx���"�v��˦iS;#R���1�g驁I
F���t��I�2#�qx���'h�=l&����Vb��	1���1�(Me�{����_�E����'���C(�� ����`f��(�YJ���e*���\�%;��B:���O���rR[\����>2�R*X�H:�J6V��E�m� 6>,pa��u!r����f���5pm��jSW���Y#�FƣQ)�����|j����|Ԧ�-��Gҍ�F�S/��h0���ًn�(�_P� ��U��r6Y�����J�H���X�����4��}A�Z?�Z�E�y֚Kh��E� �,
u8~x*#���i��ձ�X�5�!�`hJ��$�0���"ӛ��$���u,�׊��U��r���i��xc���o��.��ƷD�,W�UB�-����HGԃ64�� ah�p�1���&iS;#R@�{]��ձ�c��9V:bj�Z�� ]JdӚH1���e��� C-#Ʉ�����VA����7��_V�e�^�4���1�����Y�j`C�|���X2N0��n�����a3�����{h�)�$5đN�a3���3,v��I��a$[���_�?ڑ��H�_K�4���1�����Y�j`C�|���X2N0��n����a$8���_�?ڑJ�H�)�o<�+���~�eq5x^�-i�I�<Eɷ�O���!�c��y0�?��!vG.Si=�՟��I�G՘�&O|��L����ۦ�?�l&Mqx<�3"&=e+(Me!�e	�����=����g�D�����K�\����&���"c�RVP�YBk.c�Cv{������!�&b�@ $퐘�� ��7�̈�YGJ�Ue+)U�&��H�)�'��
}�m��qd�%��4�+��ߌUi3Iϛ�n���u�cW�S0�i�	?�=���}B����?�R�J�Q�+�~0���1�$����T4����v�nF�{/���qF�}i^i3H����݄�7)�w�?MLzHR7�@_K���G9}/�S���'�����H��;՟��=$}ox���Hia$s�⛴<	��#{@�V���g�I�@����I�~��p�&��YH	Ys�S���_F���E �C3��'l�� $�p���&dD��:VR�(qYJ��5�2F�N�8��p�S�Co����ڎ�.�lװ�.�h�XH���V�#з���n�+��@��B���2�w{��\xo�S?H6~�w������S04�$�86a7Qb/�I�p�Uj"܍��$�0�lt��ܣM��P԰i^J�D[�^iV~�r�qw�iQ_#O����<J��Z\@Ң���T.�FG%�z�3x��-d���ԆZ+�d�r�qw�z��jv>o�P��V��1ƈ�C��He ���B`z8LL�2"Ue+)U�8��VP�˙#d�p�GS�|)�Z���C
O.+J�|���' q��&i $�w��L�y�r0���ل�DQ���$@/�.)c����Q�m�A�����Ƌ��A���iV�K�*+̻����RطaZM&~Zx~,]Hp��46�*(�_PiQ^f�&�-i�W��q�K��ZM&~Zm���A���i[����e� ��!M�x����X���>�BY�2���YL�Hn�H��;՟��=7�� /��B�$���pq���6	g4�!��-��_��XoI��Hz�7�1���_K�i #	!ů�����G9NrF7 Xn�0"���
n@�����
a8�0)� O�����!N��V&}��L�'�DǬ��e	��5�1�&�Wpl �.��#E?ׁs?)�v�LOG	�@I��fDJ���e*�����Ys$l����w�>�T6��aH4�Y�f��c�Pw
�Ԇ���.+��$\VPqf{wڴ�}�lQ����4�Afg�agL�}��PiQ^a�%J�f�fG��|j���]������)�7�����=5��P�����)�����Jl=�5�SPo�,zj%3�H�~1��"�E�	"}.1UZ��#e�	?�+1ȴ��X�����4��}B@h��kQ�W�υ��qu,T]��D+�*��L�E�q����4��}B@��R���3��G�|n.��J��wU�J�"̈́���J����a7Qo��T]����jX�<���jd�V|� ��_Pm�c���R���3�fx+I�E~Zm���G��w0��]���_��f�e3�5"�	]\`/0爻T���+��!�	 nS�V~����/x���I������x�%��B�t"�/������$���zE�	#�����d�!�4=V�0�Z�_�{�XoI����}/�=d�t��PY���U��1Ɖfl0	���P	;d&'��� $��3"%VQҲ�YC��Ue	���6Jw	��u;�E�|�0�]\V��/�H��	U��$Y�7pm���'�Il$�86a7Qb/�I�q���E�f�e3�5'C	#�S ����܁ԥI�a$�J@C�B�� /��/�I�2}�)�fl0�/�'������#E5��]�'�!�N�	�@I��0	3xLȉU�t��VPⲕYBk.d����p!N���j��9)�.+���+�|`Q�0�X���wYJ�RA�kaq�E��E��U�/�ƈX����z��j*ר�� 4ѷH:�J6V���{Bf\��v+|d��(���������ZL�.�\X)'�)�*��,��L�ʔ܅ł�ǂ�)��i�$�0RLZCh�>,pH~,]H�ƒ�E�1�Y��Ȃ@#|�T�"償��	"Ӛ��W���<w��l�x��Z��0eg?$�i���Wu�Y�l�f�ԟ���K�)%i1XI�`�b�V�e�^����ξ�`W�9j�D[�͋pQb����,.�������-ɏ�{\�K	 S�`W�9j�f�e3�5$�@ܦ0�Y���?MLzo��@_KI��i�$��}/���@Y�,��G� z��R��XI�gܲ�8�Nk�N�a7yz��R)��S���-��_�.���H�_K���H��K5��5g驁M����`@�8�Y�"����/�����>�J^p=���ҕ �������	t�$�r��L �����S2)�
fE0<���ҐALȧH�a$~/��f�N��V'�Bl&M���П����&����1�8@w���`&��� h�P�2�@I�!0	=&&o	�*������VR�(Mȇ�S�N#��>�-P��!�'�հ��@�����f� h�(^�Sc2�=���M��D�a�4�F~�/w)��H/��/�Sc2�	���q}BH�S�\[�������ֈ�.�q�LVr���W�U@�b��ǑLN@�z�&iS;#Rr�$��Lءx&v�����*NU�����l����`Sr��X���I0��ءx``R�@0���3I.��a0q���1�(qYsÄ)�����1)�v�LOG	�@I��fDJ���e*�����Ys$l����w�>�T6��aIa�a �X���&i�¬��zx:���#���=�3<@����P���'y����4��~,�뺈�q}A�E�,pp�T.�.(�w�j"ܜ?�qLN@/���ZC�	?��r���J�o����	��MO�����E�'I�����2�]X@�u�0���'����˚���̈́���A�-(�W�C����T\[;Z��+W,���W�� �� ��w�R
�Y{���G��0����$>VP�Ys�"ý&~��^9�E�(,��!�Y
�hwj"ܒ�e�)�~�p��<��]�AⴇF~0��b� iV�K��8n��Z��#oqqZuVjvzJ�,�I�`w�ЋOŋ��J���.l�j"���켳�`<�T����E��H��ߐB�/�sga,��?դ�"�gdjN�G֦Aי���܁J���H�)I
F���t��G9}/�S�������+�*�t��?�B�	 n��=$}ox���IIZ�_�!J�����S��}�0)�B�'����4����a0��	���P�	��Ӎ	��%�'���YC��YGJ�YGJ�YBk.c�p�Gp���t�{]�s!�;U�����nâ�]�G'	�c�S����|E]�l)�h�A�?f��'l�� $�p���&dD��:VR�(qYJ��5�2F�N�8��p�S�Co���ۨ�j~��jG�_��ź��fȃ��D͕jX7�\^mP���MH���7]��4��fȁ�H����ZL�b���#�n�J��ga�`��
>E6,*�~ŷ�l�J��Ҟ��J��/�4�����_c�=�[q��*k�c�?��Ja��a���x�V����
mw 4K��u(��E����]�i��ԃ+�D�|��:�u4�d@Ң��Hqe�	��HpŸz*�(���#�k�鴨��v��_͋�^� ����
F�m�iQql�"���&+	?�ۦҢ���
>l�0�X�����"�o�;�"��u�� к���I�Л	��Ӎ	��	>w�=	�� ��DǬ�5�&����&��*�YC�˘�!��ʧ�ڔ�-]�\i-إ�c
4wP#��D��C(�� ����`f��(�YJ���e*���\�%;��B:���O���rR9/ҭr��RZ>�X�,$�<b�I�E�������G��T�I��O�Gz�� \Q_͍Uj"ܓ��O�A�D�.(��u���8Rj�D[�������0��@W��z��������["*px�n}zL S�g`ѣI����b�B�b�R�f�8~x��(��F��C�����Vb��	1���1�(Me�{��mS�(��Bm�tRk��2�@I�!0	=&&o	�*������VR�(Mȇ�S�N#��>�-P��!�&����K�u�X�:M��g��y����4��$�8:��&-{�"��ӻ�4cc/�`Uj"ܭQg����]����HԒ�A�	��k���!��a79��u�#��}B}�ұu ./�����+Hya�&����+H2���s��QP��J��Ҟ����Ң���*.-��U�����i1��+�h�_Pi^1U�#���ǋ�KV|l�c�?��Ja��a���x�V�`�OÌX�:M�K�
1Y4�y��D7O����r��T\V�U��������~,�+���q}A�E��,y����=���E�8ư����a���R?<�h�/�d@$yUj"���Y��b���4��}B���yZL��$�.�&����bM�s�1HRb�"�QfÁ����0V�4����V&7Bp�&=e	���`"]�J���/���"�!�N�	�@I��0	3xLȉU�t��VPⲕYBk.d����p!N���j��9)˒��۰��_HW���yv�&i������S'��uf+	�����L���	���6)B����8��5�p��5�&���P�˘�'��>s�|]����ߏ�qn��2Ɗ�1o�"�!�N�	�@I��0	3xLȉU�t��VPⲕYBk.d����p!N���j��9)#������i[��qp2�H0���6T�F��Q_�*+�i�����+I�Hp'��%39[��_�6�02�IL�sI-����&�"�E�	"}.1UZ��#lV~T�[u�[mZTW��Ic��%��*�֢-��f����u!����?�1*ZmN�R2�+wSL��԰i[�e���ZE^�"�]�ga&��,�i3H����݄�7)�w�?MLzo��@_K���IM���	a�l�i!v:o����zLvC�a�!�����_�{II-}/��,7�~��9�s�0)��w )���`Sr�t��@S	�сM�|�/�&i:.��a0n/�����L��	�1�(�YBk(Me�{���O�C˰�����E
C(�� ����`f��(�YJ���e*���\�%;��B:���O���rR�c��n��ƥ�J�̱� 6.1U��"���u�oA)�.i1XI�pl�]�E��D�M��UCK�4��Q�m�c��85�Ǎ��,W5i1XI�p��H��]cWyc����ޗѪ�E���`�k�h�4�]vn1�`ҭ3,u!���aF��f�f�O���Wk���^���;�AǇa ��"^]"͋d�hw]���i4�jXH��H��LG�Jů�M/�PiR>�%J�f�e3�5#�	�5'C	 nS�yS�����%l%Dڑt�B>�68Lh�2V��L���t#�Sc��5��~��b�!���/��;E/�y�J�J�B>�7��๯�-GT܁�)R0����7z�_��
g�N���H�_K�_0���J���`Ҹ�HÂ�9Ǖ0!�#�{���GF>jB�	#����Q�m�Yq�N0O�I0�`���L��_�H�t#�_K�=[�)x���JLp]^b����*���:��lg,��z�3=)2V�#iQOK�W5iL&n%#Ʉ����I	��9r��ʝ&iwVb��	?��!�?�a0ct&�`$���T&dDǬ���5�&���Q�Ys�S�پ�<����yF��'m��v�LOG	�@I��fDJ���e*�����Ys$l����w�>�T6��aI���=�Lr�aqvv�/�5Ha�Ƥ� ��O���c�m��l�VnO|��G����A��fj�&���S���/�}�z*�i0��t� ���vD�`W�r�7���$ ŭ+{\%J�I�=�݃Ȼ	 \QF-K	 \R� �&���6D+1��1n�i�	?�H�
74o�ٲ iR7�%J�=���t�//Q��}�͑J�4xJ��� к���I�!6'�Bl8��{�!6&j�&�DǬ���YI]e+(����S�Ys�;n� K�XNY��Ɵ��K1�$��M�o�&�`$Ǝb�	1��DǬ��e+(�YBk(Me�P�˘� ;�:����������x!O��g�	�d�	k	�1�(=��������P�˘�����q�"v3�CBv� ����_�߀"�!�N�	�@I��0	3xLȉU�t��VPⲕYBk.d����p!N���j��9)#��E��5۰�v�P5�� E#]v�m!��i3Hqj�_�	L����DG0��P	;d&'��� $��3"%VQҲ�YC��Ue	���6Jw	��u;�E�|�0��?ZW5i3I��5� v�X�=�MD�`&i�&|�ZC�U+J�},p�`�*]B@㖤X�k�/Mύ��i��|��r�T�J��R���T���9볽��[J�}k�X�^j�XI�,$��J�̾�q�G����+H`�H��H~����^��J�-�vu�9jB�Mz���Z���G1�	!�ҭpz��#���V>p�	��>s�Bl&	�2"c�P��YO]e	���˘�'��3�4��XE����� d�b�@ $퐘�� ��7�̈�YGJ�Ue+)U�&��H�)�'��
}�m��I�ϐ��+���&i%s2S+sI�a'�@ɷ��"x((�6uǛ;��-K��cXI�i���r^7߀@ɷ��%�]��F�i +��`iV�f�O��L\o�� d��H�u4�ۼJ}A�bx((�Pb۟-�s�/�Ң�=���V�4�)���:I�2-"mK��j����J�J��"儐�\؁�q��w�a+�����iR��+�k����S����B��$�p�&��YHaYs�@G`�2ƋH��1|g�xP�2�@I�!0	=&&o	�*������VR�(Mȇ�S�N#��>�-P��!Ґ�H���$��i�@�I�l}��l��|?�	�K	 R�'��a�V�4�m#��>���L��!�ϼ}�1�rS0�i1�$�0������U�� �҄w����>�-�� ɴ�Ei�$���p��"��D*�c�o胍K��D[���'�`Ҹ}��"�gdjA���M��F��W��s�����8���Z�� �.-GP���w�Õ�;�I�ϼ
W��s�n>���%�a+�$I���"����ѫI�Hauf+	��>�p�&=e	���`"����cE?��!�G�'�!�N�	�@I��0	3xLȉU�t��VPⲕYBk.d����p!N���j��9)R>��5⾴���c�@�P!�G��$�)�_ZC׉@԰ ��������c�@�ZL�#��r��O	jf��l<�MA����nC�����ju<%��A����)t���6�01"S �!�G־����D�L��ea'ᄶz��O�Ѵ�n����q�D[��F
ҭ�{E�û1�A�;ۦ�2��/nl�%0�{�Ok�����aqL�� ԰iV��Q�D<V����$�H��]f��oK��;^�Mj"���-�NE}iQM�M"�����"�����5
���]��%R�fsH�`��خ��M����T�)��%�g��S�9X4���^��V����&�[�����@�/�_�S�_ZW�Ej"ܬ�,���H��������هQb/�I�q���E�f���O����7 ��� I�H�) �5,p_��z� �b�D}mr\k~G�@԰��:���i�$���4x5����6�P\@(���>��m�;
�(�m�"��n��[h�m�{v*A���V�4�)���L��:Ir��ʘ���ox���I+a*&ԚLt#�Sc�Ǝ3%j~��Huy�z+�J�h�H�c�Z����tS�Ǜ��t��}/���)xc͊T�V:����/�~�j8j��QJ��8�^��R�0S>jt�&G��]$>0����~X4�����
�0���Nq�LzH���}.�фϚ���H�)���u�vDb�S��RA�%D�.�`m�>���3u������� ���=��x�V�h1Ўw�~�)0l�#iQOK�W5iL&n%#Ʉ����I	��9r��ʝ&i��1XL���l&M�!6��A�?f2"c�Qme	����YH|���a�G;�9T);R���F�F���u����2�@I�!0	=&&o	�*������VR�(Mȇ�S�N#��>�-P��!�!���E�4�i�԰�]�'߁��@���+��V�4�2������Jg�� ~N<��t��?�	L�t ~LĉL��H`�OÇ�݂]DQ��� 
g��_X7�,�8-D[�qY��]�0��%����9��Kԋ6s�3}�%���%��q ��դY�����a/`�D���(����ӳ����D[��g=�}�E3���ZKV~�,e�J��������W�>*�D[�W,$����R����`W�_�ʭD[�Qa'�3gK��W�5�_~pw*�n\3H������H�?L�0y�������H��4��@��
jt�&@��y��!���V&?<c  ~n Є��	�h���)�\ǿ�Q�����#��He ���B`z8LL�2"Ue+)U�8��VP�˙#d�p�GS�|)�Z���C
H|Qأmv�~
����!��]Ű���4�+	?-�'I{h����v*.)c�W楇U-@X����D[���H��H]͏� �ّZL�,�vF��a$}jd:�-�
n@�R��a$r�*L�@��1XL�~��4Lz�V\ǰ�
n�2F���Eg��6�	��C(�� ����`f��(�YJ���e*���\�%;��B:���O���rR\��oijXH��e. i\դ� �o(ҷ-54�_PiQ-%i?�؀�Q�n>o��_PiQ-%i3I�!�|F����KFj=Ĵ��A��N���=&�D��rJ�w��[	��7l}��}�\_�L��H�a'ၨ�/�%�a7Qb/�4�MW����`ѧ�_Z"ܒ���d�vX���դ\����7c���r�+{J���gv>�mj"���S9Y���}(���0�Yݏ�R?XI�4����݄���,�U�� �ք�Z"ܭC����E޿د2��wq8�*�i2��%�J��k�����D<�!�`V�a�3x�c����zi�$�8��!�em�v�Q�ךE���Ԏ�&|Ԑ�	!���#� C	:}E�f��	���!��������lM�?�L$�r�%,7i\����S����jN{	!ĺ�&�5:E+	!��t��z������A�䲃p<���H5���S#D�T� C��D�~b�ZC(�� ����`f��(�YJ���e*���\�%;��B:���O���rRb�V�b/�_����5,$�om*+�3�p�$mI�h�w�Z�I�E���m��#�]3Hr�O�#vA�
1��U���wj"��s� �	�߁,a7[�A�7��0Y�7�)S;#R)XJ��y�� a�ZA�	�����IM���	a�l�4����h�ܔ��:if�6��/��0�r�L8]Z�<� �����c���� E��
4dFB��'l�� $�p���&dD��:VR�(qYJ��5�2F�N�8��p�S�Co���){�"�[$(����$虞�H�ؠ
k���O�o��?n�@�Dfʅu�v}�\r �+���}�ԛ����x��95����#$A��=�=-�ZL�cH��&�H�r��4R��Mx#�0�!�����=�Ʈ1bx�7y�����Jda�G�	?�6���M�MK}-����/�=N1��V�-�^�I�)�E-��G��X/��D��f�'����Q����=�dx^5����A�縘��=�����j%j$ʕE�>��v*�#���]���Ң��,v�jE����%�9�%��'>��ρ.d��3�� g�rs�TNi��k;���]�k�_Ph�GY�9�����~��m�l�^^�H�a��]���wL���%���E#�F�,p���'��_��iQF"���p���a�����sRh3��6v*(�_Pk�!�F�2��~�c��E�8Q۬��4NA�G��kv�o�/�|^�k�&�ZC�	?�5�h�XK�
4E����`����}�%}��}��j2�E�t�&�pm)����Tv��u���\T����ⵄ�<Oi=���r�YzҢ���#���#��Z�2V@޴��+"�QZC�8\�����qs֕k�����8�_������ȑs ��l8v�c=Cr��G�pw+Htg�O~�S.zҭq0��׃u�+�`V�A�5�F�KA_��;؟Ã�ZC�8Q���50��*�,-x7Yq���qiS"K�cPܣ��8;���g1�18�r�]�^�+ۤ9�A�ԅ&�+H2��g�I���ߖ����u�+�7N5!�
o\�k�
����&/�԰}�̾���IZE�8�Z��ja��ZU����?���ҭ��UZLVq��c�#Ĥ���n�{mv3������e �z��� ��ޭ�O������F�\��Z�ȀH���+��"��@B��f�3	?�'��R? ��|�i^3�U��rN�8�����3�a5a4HYH|����)㱕����<t����b� iV�K��8n��Z��.��8�����-�N�Q�'af�gaǤ�&�	?�z��/�`E �)ԹV�n6v�y�H��U��s+�"�gdjLV��#_y�j8��ҍ���e�dC��a�HP�9Až�m�ڴ�+	]b���� ��>���xY�,�,DX헂�b�.�m
IyZE�	 nS�iq�N|0��~.TN|\����s����V'�֧�#>o=V��#>e0!�^�}.�4����V&7Bp�&=e	���`"]��1ƈ�)3��'l�� $�p���&dD��:VR�(qYJ��5�2F�N�8��p�S�Co�����[��TW*Åi3H�7)�#�ey�:0���݄�9�E|���O��ʛ��e��sY����	ZE�1�ń�<M4�6c�������a��4��[د2懹bXY��w���B"���ǖË��A�w�e���7�
T��1�Xqu�4��,��Ң���J�`�}]F��v�٩���nX�u��Y�%?��3a��O��;��V�o��tCJ�gHtf<s.�5��E�ڴ�x��W:H��Pa��n|�j/�4��1�`R�q��Q��_PiQ^cx��I�f?3.�s��Sm�J��^`�!�p3�Y�ia��n|��ڴ�x��W:L�,�vF����jHů�q�ܦ��&-!��K�s�ߛDv
nJG���s��2����Sx� S�9b�9�o�q��nSp�����jn@�����
`
t�&7�4���1XL���� �('�&�` ���L���a3"&=e -e	����YLz˘�|�����v�����>���4��݆��v�LOG	�@I��fDJ���e*�����Ys$l����w�>�T6��aI�>x<d(�ZL�@���Q)�a�M&~=L%�h�?�N�|Q���+�/��E��1�*-�@�h�Rf���c=d�l��Q�A��H3c��-����n>E�{�A`?��e��,t��c��a�6�(�L��|h�i,t{�Ʊi�[���VD+q�ƋV��Ci�H2q]kq�,0��Y4�{[��c��e�w3�n9;	 v���ZL�/��E�t��\A�v�,8ԋ6:,��M�ZT_`��*�WZ�,@g�PY�;�~YF�íx�e���`�=;	!GP�ּ�3V�J�C�͋+��x�l<�RդR���`ŕ�E<b,wL�
�nc���+��x���frjZ��Lt~`#/ 4M��`�䰳����e,
�X	��E�N%���Y�H�
:�
�X	�m����+7�ۦP�\��uۦP�� R�a�(�7�"x�`ݠz3��DYd�4���^�8ԏ�:��>E<l�8>j�?��t�g���)�d@"�+I�H5�q:���jO�:/���ybی�Sօ�����Pc���Z�+�
>2R�5V��EX6 |��T�u���I�
?$�0�դ� �����`+�@ i��hɊ� 4��w��"yI�b֏֕S)���jL�nb����L�[ۄz��f�e3�5"鄮��C�9
6"��Ƌ�a=��Q�H`����5��N���Hjk9j
t�!����n09�`P�)�Ё��l������Xo��|�B���L %���9
6)��a$=V�f���V-W���&È@ә�	��	1��Oq�&��Lȉ�YBk(qYG�e	�����=����ӷ~i&���c�LCg��Fa0Kza0�XW��BfDLz�VP��J�(Me �˘�"��>r�mݩ}�;���DA�LŤ2�@I�!0	=&&o	�*������VR�(Mȇ�S�N#��>�-P��!�!��iV���Fz�^�4_�'aÅ&�Ѩ4���*���vû�ZL��:���4Z�����)�~i�$�05�h��	{���^�4Z�Q��a'��8{�B��i�E��`|�-D[�� �d;�Aډ���t�ݎHtd>7c��x����zC�!{�&�a��	��>��.���^��	��q-��}@MI��_}@M��{�&���d/���&�c��	��PE�f�e3�5&+	]\`/3w�yk��6�L�:�դy0��]!I�߭ٸ��9���u�N��h0�9�d)��s�5����&u[��|���$�r�J5q��h�Ʀ�	�V��_�L�.��a0z.a0C�	��'XLȉ�YC��YBk(Me�\ǰ��p�SOwk�ȳvN���#E�Ť2�@I�!0	=&&o	�*������VR�(Mȇ�S�N#��>�-P��!�!��n>E�i\|+w�����%$o���$F�5ۢ7�l7M����IL�\�8�I�n���%dJ��/�_E�X`���nI�'*�"7a"Hi`����~=��rË��|��>��.���%���7-z�&���`��8����Ma��t��A�Q��i���.�4��$�7M���a7Q���U�n�,A�����nec+/��V��uٮ+q���"�#E��X��&iS;#RG0����7z@��/,&��<�M�.���Hun9��n�x���$a$>�~�H]���M���x�%��C�zO���	a�l�i:�G:z/q�����rRBlt!�>��X�>u&;	!���f�����I�a6&uP�	��2a0C�	��'XME���&���P��-��5�&���Qme�{��>�h;_nG���{�4��vdf< �G��bNDǬ�>��=܏�`#�#E8��5�~R@ $퐘�� ��7�̈�YGJ�Ue+)U�&��H�)�'��
}�m�J�:G�$���4�j�f��q�A����ף�{�#��L�Rg��f��}��k��=��D�~��_���M���7M�O���@]vha��nI��5,V��^Z���ZA������G�^��&�-3���U�԰}�0-U��s+�a'�#�0��.��?�M��*���]B�5gkQ�n+��xG�^m�n>n�W� �`�t��ҷ"�15i3H�a'��n�J6�wRB�ˈ2寭��3��b����,���E&�Nв����_�|O)X��b�+\w>w��\=i3H����9���0����1ya5V���n�t�����n09�`��H5�������:��lQ ��a,7��uz��(�joI�t"<7Xo�N��c����3Hy����A	��!��L�&dDǬ���YBk(Me�\ǰ����{�)E��k1�!B>���Bl&_��0������YLz˘�r?��!�v�Ɗ|� �'�!�N�	�@I��0	3xLȉU�t��VPⲕYBk.d����p!N���j��9)#��J�ƥ�J�̱��a q��&�4SL���U���j�f�Y�u����c������h�A�k��v����Jd�L���Pv��aqp4F��5�@;a�zj%3њLV~2WuF"��� �����Pj�\K�A�r-D[���./�G9����J�f�"̈́��
,%�"���c�WX.2X�i���j"܏T��K7+H��O��9 퇑��mZTW���#-D[�X��9 SCn�F��4��3�ZC�!�
hm�&�ҭ5����q��1�H?��F0b|}��ic0�#�b���f�e3�5!�	 nS�V~�����ox���I����_K�.�S_/�_/��
n@�z����u'�����H��;՟��=$}ox���IIZ�_�!J���H�HR��XI)N�;	��M��>�$��q�����ܧ�#Ʉ���i3Hw�Y��`!��(G�&�` �Bl&<�̈������YC��YC�˘�J��k��7�%�i]F��p�� �w����P	;d&'��� $��3"%VQҲ�YC��Ue	���6Jw	��u;�E�|�0���]��K�A����԰iV��85,$1U��F���N�/h���[�n��&iH�{��6��~pjr �>��l<�MD�W1�h��859 Us\��G��S#<�~2WuF"��� ��b�U��r6\������a/`�DQ���c��X�nG�d�w)���l�wp���$YH	Ys����f�OÅ��}@Q���+�,p4��`�nG��f������@C��w�M�e�~o�N�0������H��O��9 퇑��mZTW���#-D[�X��9 SCn�F��4��3�ZC�!�
hm�&�ҭ5����q��1�H?��F0b|}��ic0�#�b���,�vF���&@q���Fq���6G:��5��|��|��	)pF���L�_/���%M�RC!H`��j���5N�a$s��S�Sr�*N{	#E]��h �)�B�&iWVb��	>w�=	��&П���*�YC�˘�KW}��-�����&��)���l�wt�P	;d&'��� $��3"%VQҲ�YC��Ue	���6Jw	��u;�E�|�0�{e�_�LSA ��?�D��yY�����<�P�ʫ�����/X<�_'�9��V`�	!�������[O�v"_�)�L�1���(��e�D�U{c;:d(9� ~�+�o��9��Zd����6�l8j����,�P��L$��U")*��0�	#D���]�<�V�@d20�����DӶьȯ�9��/�.�@\,�6>�p1ŭ��V-���Rc�侗�"۰2�e"����Qu��.Yr��u,4M����V`�a$.��Q�D<U��� 4p!pz ��Z&s����:I��M�E��0��%m����J�1�j&s����W�GY�V_��X�!�_��Q'{����I�G�\��}�K�F'"�H_'�P��$���E��4����+!�>B�D>Q3��X���N�@�F�1�L���,�0ݲ�I�II��L��V�����6y�@E
C(�� ����`f��(�YJ���e*���\�%;��B:���O���rRhcv�a�k�a 4j��F@�F��;��C�a��f��6y�C�<��kaq����I�q#	����U�["�õ17 Hz��We��r�R��o�@����i�$��I���Ë��1�ˌ�3<[���Z5��v�	�j"ܺ��J����P��;B9P�R봾eO@̠�3�5���f�ⴙ�YL�HÂ���1��o��.�I0�Cg��D,7�,7�N�i1�IU�����Vb��	1�	�h���&��=��w�71Ƌ��	���P	;d&'��� $��3"%VQҲ�YC��Ue	���6Jw	��u;�E�|�0�\�JvqF"��Nݑ�G8��F��T�&i1����%3+� �a'��	���}A�oRó��G Hz��We��sFVc��Z�~(~+I�E���ԅ&G9O{c��܁��\�s��
{�u=S��#���V'��'��6����B?!?�&=eU�&���Ys�	j�ҋ�f�ǀ�&���{�������[YA�e+.c�`���B���F�����f-!�N�	�@I��0	3xLȉU�t��VPⲕYBk.d����p!N���j��9)W�n>�	�D�&i=b/�Do����4��~����o��>q��-�f�f<F�$Ai�x�,'��
E�c�����e�m�"�1��j�e�m�"�1�Xp}�����֑a��8��Y}@[EkI�A�	?�+�sC}���]q���/��u����c�E�����h���?���+q� �+I�E���Ԑ�	�ۦP�`"�q��O�	#�"�q�� E�����q�Y��`%��b�l&o�����������P��B�1�=�����1Ƌy��&b�@ $퐘�� ��7�̈�YGJ�Ue+)U�&��H�)�'��
}�m�8��iV����,$��݁�ZL�<���w	h�����!��O�KF�n�dQ���Ң����ʪ�E���e3�5$ �H�o=��=���=폺��f��uf+	���x�P�	��s�~xh������*�YH|���a�w�iE˳+1�&#�s	�� BDLz�8VP��-���a4;�Jh?���cEs�G8E
C(�� ����`f��(�YJ���e*���\�%;��B:���O���rRK��J�u��n���ҭ3h��Э&i�>ds��u7��N\j%2��E~FJ�(�_Pi]K����*���U��s+ư���0���1�U��u/�j/�4�G��V�-ϯ4�6~]A����iԿ��p���s�G9���21h��g'`ҭpz�\����I�n�W�N���˅��4�L�:��f�e3�5$�n|��K9�`�Hr�Hzl7K�`�1j聉����PP�$c���1�IU����~�Y��`$��6&�Bl&O��OEBl&�M��A6��Q1�(�YBk(����Q�YBk(����P��=��f�)�gk��Z�Pr#�ݨ�1]�ُ/���NDǬ�=e�{�|݀�������P	;d&'��� $��3"%VQҲ�YC��Ue	���6Jw	��u;�E�|�0�n�j�������l��5��&8���������N#��E`W�(X���Jdg�O�~}8���uF"��J�k��*�nFج$��V8{a/q ��G����̾��"۰hǁU��rc�g���6�M1"��pT/���"͟m��F�ga���}���8�!�4�Ei�$�(X�턮d�v�:�QN�q����,�TM�E�1���iW�ҳ��RP�͗���"�gdjO��}�J���)��
6�]�J�=9V���-+�q_K-������J�=9�%�f�[�1XL�0~x�>�&�`!I��'�DǬ��e	�����atPvS���P����~R@ $퐘�� ��7�̈�YGJ�Ue+)U�&��H�)�'��
}�m����v"	")`S��{]�jXH��7듰�0��b���P��iQF"��k�3,��.��x�V�4������A�����D�a���5��M��p�)G� �6Jgt��h�l��/�M&~<�.�*��{]�Y�P��j����b�����r�r�Eu�v��89�@̲����V�������6���,�������P� ��ڡu���rp0`�qv��@���x�>c�@��и��I��E�}o��>����~��M�E��D�B�88y*�nq�a'��Ȥŕ�E��(�Q�V��b.}F�	Ɨ��c���n7��~o��o��ԙ�YL�H��H���q�����#{���Hp�o��_�/@��4��Vb��	>w�=	��#!6.|�΄̈���yVP��-��5���\ǰ�Z��R���i;9���Q)�v�LOG	�@I��fDJ���e*�����Ys$l����w�>�T6��aHt#a} \4��ȼ�B�|F��!���Ki� �� k�}�.V�4�[������}����_G����ޏ���D�M�H2������En�v��J�X�
s �v��"H/�4��03Z��+N�����`�1�4�
v�}i]K���i?���X4��z�_J��L$�7e�x5�����4����(�+��,�03Z��+#�aq�/�4�B��+	?��ޏ���IKq�n�L���`Ҽb�}�3Z��+#�aq�/�4�B���ư��V�q�EkJ���xr�i�I�_�n|�*԰��iV��W�ZL�,�vF��a+���n�w�^XMU�y0��]!M����n0���,�.�{H�c���X��r���X"��a�����A��S�,7�I1Ё�� ���,����XoI�G�՘�&O�a0gU	��	=	��#!6>p�	��m	�1�(�YBk(Me	���e	����YBk(Me+.c�Mn��A���t��-�������`������Ew��!�N�	�@I��0	3xLȉU�t��VPⲕYBk.d����p!N���j��9)4����ȇ�+��uߗ�#E]��F�x�����mu�zzv�^�W�J������ZL�(�Y��`$� �dG�&�`!��(G�'�DǬ���5���˘�|��%�.]���� f"�!�N�	�@I��0	3xLȉU�t��VPⲕYBk.d����p!N���j��9)?�) ]�,plPQd�{qJ�f�&iR~�)��q����G�H�c�}�{��F����_�j=�����;���^���IL�f���O�E6J��;���f��X4���j"ܒy`��״�2�H2����}��k����F��+��L��]�}A�n�86((�S��Z��2�&~�^�㾆u�/X���V�Yc�b��%;�,�U��}C�Q�V2�K���9w�.;��TQ���H��g�!��/�~�z*�/�I��L8{�w���l�J�宻5@E��r�f�.�.��I+. h��ZC	��i��Q���A�EV���%J�8�I�`k�qu}��W�J�8��� �AU��r���OÇ�C%wQ��dC����Ҳ3�,�0PUj"ܒ�a'�'r����n�:Ml,�*/�_PiQ�H}��԰iQ}���V�-̬�BC���u,�H���Jw�j�f�ea'�X\i��)ƥ�
K�F�J@S�Ѩn~i�%��V�4�)���#�J��y�� ]��UiL&�=�簒{�����&M'=��3�����L��Vb��	3L&�`$��&�`$�P�	��2a0C�	��'XN؉�YC��YBk(Me	��5�[YBk(Me	���˘�!��|)����J���Q����Owk��,��Y�:��؆�a0�Oل�������P��c�\ǻ������i	�� �"�!�N�	�@I��0	3xLȉU�t��VPⲕYBk.d����p!N���j��9)�*�1~���&i�}��A�縚 ��?F�:�!���
O�)����q4A�=����mu����/�RY)�Te ���(j`_�Mlg�K=�%����>�r����E"R��%���%���S�#�����	{F&�Q�E>m3�T4�Z��#a��x>jV�1N�π/)ga ]��Mj"܍���eU�菚��5g���r�����w�����3X���^��3���
O�7M��*���|��>j�?XI�	�K�
17M��+u"i������E�i1h�D�a-3���v�95�u���iD�nFج�L�:���;	 f�}�<�CJ*A�.�1Mo�bYπ"�)B��@��ԭ ��O�A��G���x��6�4�L��>j�D[�[������k��약���,pK��k��2��N�	E��r�-�/�]�԰�~Ƥ�&+/)!F�뱻	 �-��S=a$�)l���ф�<F�'��6a?zE�.r��4v�D�_�e�c��j��f��`�r5�&��6�Y�j�|4]&i�$�.�w�w��J�m;B�ˈ28�1X����Zf)�io�PiQF��;�	R��6~]A�!����e �d����юH�c��c���_����F-#l�R�뉥n�������}BIZL�,�vF��a+���n�w�^XMU�y0���a$=6��Cx�%�R@F:i�ޒ1Ўu����$���zL�.��a0{�a0c~a0xπF2#�a0FB����&���PⲄ�R�P��-���`"[��4yݯ���v4Q����xAЏ���4�	���~�'�DǬ�>���S��=܏�o��|݀=2ƈ��K��h)�v�LOG	�@I��fDJ���e*�����Ys$l����w�>�T6��aH�cȃ���\E���Ӱqȵ��_99V�H��ю�;u��Vz�Q��J;u��VJ�Q��)�j���������'�8���w���>n��13����Y�.��=������;���|���tL���{S�c��v��y�3��Y�^��9lǖ�ڔ<l��ø;��/�Q=f9�'���1�/q��zܽ͢��GA����k$L��g���h�/�Q�f���^a�^�?���E�{�"�s1�3��͢�F��3��Y�[���(�3A����R��g��-�������{�5ُ){����m��������d��zs���=f�z�,�4�d+R���,���&���%�pw/R%��m,�2��v�D�Y��?���q�q��%�`�\��>FcY"c���?���q�q��%��m,��2�험�=�g����5�=C����0�A��y�Z�Ã�����X�Ѥ:K�m,f��ؠ����绌���5ƱǣIk.9�iq�1�q�q谓����6�֐��..���gIb.}K�������wm����%��1�Y;R��<�X�6�֐�-����A�3�X��X�Ѥ:�^�d.��E��8=c�k�c�F����yq�1�q�q谓�<���4]!I�\4]!��"Β݄{'��r�L���,�9d�J$3<�9c�ۯZG�cˎa�k�c�E����mרa��
L2���9t�@�  u�>��w��ȏ��>,]�i�n���מ��_2Wn���

�(�Gϵi���i��X� sF6�Q_�&�V� �g� �"��
���Hn�{��^�Ѿ�dW��D�!��9�_(����Y+I�Om՘�&L�	��	<g�#�	��#!3"&=e+(Me -e	���˘�!��|U-�qё���x	'��p�&=e1�.c�|C��8
���#}�He ���B`z8LL�2"Ue+)U�8��VP�˙#d�p�GS�|)�Z���C
HD��o���z�I�HF��%33I��O�G����MG���o�1�8u��Z��#��1�E���B����ųŁy[��i,"jH�:(��njf97{HS,F��#����x��L�!��i<J����`x�H4�0�����rn���[���#p��V��c�7�#sS1�y��B�o�.���0<U����������<��'�@�غ"#p��V�9��?x��L�!��i�"7i�t:{����X�MG���$�����`�y����������ga�E&�>>�@��� W+n.��J�|��V�A���x��L�!��i7�#p��V�A��?�F�c��w��%#p��V�f�O{SS�$���}��w���qʫH2�������I(;n�A�käz�������t�,�f��c�Y���ZL�X�gO qzɭ���_�9
6�5"͎�q�{�/Y5۰� -����P���i9N7Dnqv�_���|=�դ�c��#vnzҢ�|�Dnv�95�u����ZE��K7�#�v,�zҲ�Y�/��w�>���$@[�-����|��p��i^=K|��Q�>�k���Y�`V������rk��^5����6:bDn��ƕ���B���j���x�)l�_P�"�P/�^��<U�������g�!��4���XK�&5���q��q�H��#p�rƂ��7���s�ZL�i0����\�Dn��w,���KI`X�h�
�sض���W,"�UiV~ŀ�I ��٣&+�F���ޣ��y�`?i �-iU7�	�F��&�-#})��� %��G��&iS;#RG0����7z@��/,&��<�M�.��a;ì���
c�Y�=9��ʝ!�	#})�OA����ݼ:�!K�'C	#})ڨ���_�����Ɓϋ*t��;��a0xπF2#�a0FBl&	oBfDLz�@Z�YE��&���˘�|��#���=�m��Y�:��؆�a0�XW��BDLz�s�(Me �˘�r?���;�	��_�E������P	;d&'��� $��3"%VQҲ�YC��Ue	���6Jw	��u;�E�|�0�:�����v݄�/,�>���^|� �ۺ���&�դ�!���"��q�_G�Y}�=�S5n>��x5=���>>���?�D�y�����)��q�_G�Y}���w���=���[�ݰ��Q)���b���M���7N��uٸ��* �Z��$���i`eV�f�O�q�_G�Y}�qui`]q�/�4��ۺ���&�֢-��f���i����ԋ|/=�x>�I�a'��{������.���,7���_Pi[���V�-��~�O�A�a��E��+}�եE>��`���nVGFu`%���y�O�a��Ba�a��D�+(oYs���v3a*�F��TM�ZA�������Q��,{&�Ѧ�D_PiQO�8��Q�j�����z�\V�>�����~[�*)��ÈFZ��>��)XD�	{3���:0������<V)1XCق��m�5��юH�S��괋6m�b��,�/���"�K�;�>�I��&k+"Q���a�wdC�����!фN<pD�_O�D��l;��GϿa�wdC�G�9QN���b��
�D����S�c�a�w�a `��Y��^#�
}i�J۽�[��x*"�yI�g+(8��;"�Y�&�poڴ���a'��[�ʻߖ�P���v}�D*���1N���i1kJ���*o��`g$�������8$��Ei4���K��� �`����s6�Մ�=u�7��㜦#��,�vF��a+���n�w�^XMU�y0��]$�H5Z�}7�,7��d����O����1��zn0�s����1�jzn0�sH�a$:�e��Yf��7OM���� ���R�I/q�Y��5�o�cq��������-K>��J�J��"��ۏ�������g� B�H1���f���@��c��Y�8���@��sI�c��q�Y��5�o���,�oI�a$8�^ d�`��I�E�՘�&�M��K�?f�"c�Qme	��=e�{��7C��K�+��� �`����s6�2�@I�!0	=&&o	�*������VR�(Mȇ�S�N#��>�-P��!�!��>%�0X��`�(Q$[��
$�n��kR�Q�J��C��J�|n������@�i��B��{X�����E�	�H2�I݆k��Q�э�w厰�ˋY
����m�Ӥ2��S[��f_L����aFѩ3H�c�����qk!E"ͅ+[5�c0b��<�F8:��,JI���
$�n�N�"��C�	�x��O����~+XO��mH�a2�ʞ��lYMm"����?\�2[8�Ŕ�)�'A���q-�/�ӚE�	�g+-�ز��E�	��;��!d�������z�e���St�_��N�M|�>�	g,YKg�YMґ~�e�0���%�e5���n�-�/�Yn۰iV�`��Y	|�����=�HCR�~YB�Hu���3I����8�f��0�ݻqU��{���� �e�x?������37|K`��0�bP�H�7�������@�(�-�7%'�t�A�n��x���u[���<	����f�D��-���k��D3��1���eߖ:�.-d(�����0�c,a�ġD�l��(�-�ҡ;N���7��1Ml�����,.�7x�i������{I	�vnV�4���1XL��	���~�'�DǬ���YLz˘�#�� n�������!�"�!�N�	�@I��0	3xLȉU�t��VPⲕYBk.d����p!N���j��9)?�) 
w8�. i\դ�&��q�[���<���jX�Lո�{������{��#����{P;aj05���5(���j5�~�����l��9�w���԰iQ��E�%V/-{K*���$�7e�x5����u��|�*�^_PiQN����j"ܬ��n���G�Sޏ�8iQ_�����Uj"ܬ��I��Lt{�w���l�J��/�4��qc��-�ӣ�~�]F�2�Ԑ���E&�����iV��u[��W���XaqݘJ��4���cȉI��"�]�^����ܪ�E���~�c�) q��x>
�D[�Y����Q�F��t{	jѵ�h�\��[\�c�W�v.�Q�h�aäz�T/��`�:G�����8��]���B�&iS;#RG0����7z@��/,&��<�M�.�|�Hun�,���9���Y����zs���-i70�[�|������?��R�F��L��Vb��	1�&�`$�� �T��M��IǇ�3Y	��#!?�Lz�-��5����&����&��k.c�`��"~;��G�k��?��Y�:��؆�a0�Oل�������P��c�\ǻ��������� o��He ���B`z8LL�2"Ue+)U�8��VP�˙#d�p�GS�|)�Z���C
CH���@���4c����,pa5i3I�@��L���z?���k��Gl5��b�zj=��h���E#Q��Jde�!ф���lǼst�>]���`Ң���rI������ZE~��z?�eu��|me$�-l�x8��Q�Wj�O�G�g��.��?�M��*/�G�U��r�f�O�[
6)0l���6���sω�{`��ĠjX(�H�nNX/���NÏN5&ilf�lRL�t������&{�A����yUT!3��Do��4���7�u,=��(߿�9���ZA����g��<���/m�ȶ�$	k:�e���������[7�;�x�V�D/�}A�x��~����y��|�ۦ�m+w̾��U��s�t`�z�^	u�	�
�����dC�� ��`7���@Ud�}A�[����H�a'�"��p��ux�eԋ[
6�,3�PĔ��Σ["�Q�lt`�R-l(�;(��`��j�a)%�j۶D$sn��7�n|r�Y�/+I�C�	?���]�V\@ѐ/-}o��ZG#��S���F�Ң�+\wf�i3H����9���0����1ya5V���n�t�F@�t��u�����%��I���9����y��	j��	~�'=��7�KP9�'_��]&in��a0�s�L�a0c8M��I�M��I��6d&���YE�e	����YBk(Me	��5�[Ys�T5;�)����%�ނ�o;qڣ�ߵ����K��h!6/���O艏YN}e	��=e�{������2)F�xπF3w����P	;d&'��� $��3"%VQҲ�YC��Ue	���6Jw	��u;�E�|�0�:�i[�b==;E�`_P��u%d@ҷ-3��+H2����f�Ǭ�ǀ
�ˈ0�݆�A��IM����x?��Rȏ5�ZL���}�q~��MD�y��1�����-�Q)�<�h0��Ű����԰q*�n}n6~>jV:=��6�Z�zu,$�$�Q�>�k��Q�iф����a/q�����6��K�:�+q��E���GQu�4����IP����]w݀U%�E�7����aw�Gϰ԰�եDRJ�i0���б��"ǥ��z�૭K�:�D�nV�"Muc�ƻ+I�G�	?���]󺒿�Nв����9jLV-���iV��u[��TQ�k���T�&iS;#RG0����7z@��/,&��@FF2s�K�y0��]!�����n09�`Ќ���8��x�C�a�!�	!պ^�7���cq�77�-B;����Z�)
L$�V�ӟY�����|	�� ���RJ�J��$�B���!�l�ُ!�����7Ho���y	��l��)!6:�XoHSc��ߒ�9�I�a$8�^ d�`��I�@����I�a6d'�DǬ��e	���˘�!��|2��ߵ����K��h!6/���O艏YN}e	��=e�{���������~.M���P�2�@I�!0	=&&o	�*������VR�(Mȇ�S�N#��>�-P��!�'��r�m�
1���4�R�C^�&i��ɳ���e�3��8���S�"����e�3��v,��(�_P��E|q�`$x*�nF�+	?=l&�"�E��k��iƥ���R�Z��0�i4�I�]E�St�xiV�V�Y���5���A�K�|���i[����u��"�gdjC	~.M���%���]]Y��` ���L���a?�&=e�P��c�\ǰ���t>n� ���P�2�@I�!0	=&&o	�*������VR�(Mȇ�S�N#��>�-P��!� й�J��S��������ϰ/�4d`f�&i����7=�|�z���~nj=���sP{�n���
0875�D�N���$�8:��\��Zg��T.����a5`B"ܜ!�e1�.g�4>n�$�|�z���~n�^��V�,pK����S=�݅��1>֢-�9��zK���b��)�����
O�jL�K`�B׶a"{�V�g���Hi`�XO��ф�<G���
r�Y��>t��咳��֘pC���`��+9`؇�#�Hi`��+0.,i�>t��0a'�'x���-3i�t�>�8�M��-U��r6XI�[���B��qu���vv�!`\A��Z��#c+��ZL�,�vF��a+���n�w�^XMU���n�lt]���-H�a$:�K�s�~�X�,�s�K=9��x���I��>����[�L�����)_����&i��a0c8M��I�a6'��6&�ضLo�j(���[YBk(qYBk(Me	��5�[YC�˘�!��@ʆ���%����7���<�߬ǀ�d�XM�` ��a0N��	���~�'���YCe�P��YE��&����1�M9Gf�����f�7nA�7`)1Ɗ�O٤2�@I�!0	=&&o	��Ue+)U�8��VP�˙#e�I�Ҡ��X4�M?��>�T6��aH�um�go=2����g��Ƥ�!��OY�E���.q�~Ϗ�������G���mI���R�~`1�{c�)��I�b������c���@g���@��>1�@�;��9��<�1�B8�>�h<�1o0C�.|�|7s�%��HBX��,p@����?��.XI�KP>���R��\��-@.��4c\�^���1��,$�`#��^�jX\��%�Ԗ�d,p��I��O�Gl8^�!�4�Gּ��_��E|0[Hib��+���5n㕍��5n㕉���i�����6����5���� G��X�"<g����]��O�A<rԏ�~3�>��p4}��x�}`���RI�KP���a�F2��N���� ����H���4�H4�Tэs�{�4���>}�����.��1�8��#����O�X5��4�q��O��{t>���R?�I�s��c�������sϐ���O�Z����Z��u$ь�ŎԆV~���W����f���%�|~�W�,p=�)w�w��zG١>;�'�(�����~�� }�0q�R����9��G��i�K�ϐ��O����B����_(��V�9X��������B@h�GΑ|Ţ���vEޢv^�R���#l�W�CI�a'����`iR�^��#��\�Dk�6��L�:����g���O��S�`C���M��pu
;����:��|��7�t=�9�ŧMc� ��r�\��:hs����o{�]�#қ�P�99�f��C�	?�3999jC�~� }��h����9�����C�I�a'�,�� Gϰ����iQO��=�<F��ZH�- ӄ���.�Vv��j���V~���W����)XI���T+ч���!��O��N�9��K��0���-H�a'�39��G������!�"�	?9��	j #��jX\��%� �J���O�K�� u����A��W��w�K��3�$b�`j��+��>�g4`!���-H�a'��r�=������>B
E~s��� Gϰ԰��/�KP�"�����P!d@�����K�Q_�n9��3�$bј5n㕍��K��t>��q�q�R(����9��c����3�����,f�`>�0\�|)-XI�KP>���R�fR[�Y_^�c�4��@f>}����� ���+�m�!e}x|?�/�I�iuD��>�k��i���@�>R@�-=��r�/�&i�r@���ӿ�t."�������f��h��9���%����rr� �x/'
N�E���1�@�8� }��4}��x�}	c0,ps�9���C�H3a'������%;��x�>���R�f)*A��O���E|�q�Ŀ��r�(_Q_1)3Hm��w�c����r}) �C1�mK���,pN<�C�	?�3�99jE~� }�,ps��A������KP�0C�.|�>�$���%R��9C|�K�IRXI�K�Q_�n9�I	��g��G��H|a'�C��|�!�-H��OØ���r�c�>���4}��x�}	j X���sϐ�񄟁���ĠjX�(b���a�a-@RT�V~���W����A��c�� ����,pN<�C�	?�@�x��$�g }��h����9���s�!��a'�G<���(����#��jX�( �J���O�X5��4�q��L�r�Vb��	v�	�h�����.cߢ?��&���&b�@ $퐘�� ��7�̈�YGJ�Ue+)U�&��H�)�'��
}�m�J⴩5�,p]�/�H>Rj�$i��ZL����������GϩD��sW�S+��~0����n�]�Zj��/�H%V�-�1�I�	h�+��������!�Uj"���$�|��H<7a/`׫q�8%���׿�P������n}y�U�	�ǐ��cXG��z�~!Ij�Cqc��Y���DC�� G]ZLk��.�!�]v|��Q�>�k����YL�H��g�II�7����=��9�wQ ��E��)5	~K;Sr ��/����4�K�1XL����L�P������8��5���.c�p���|܏�k�c�B!Fk8M��B�}/�!���������(Me9��1�Bn��Q��	�����B��'l�� $�p���&dD��:VR�(qYJ��5�2F�N�8��p�S�Co���26iV�_�[~_P��6ڋ�]�}�8�!����p3V�4�K�?qj��}e�X�}=��j{��=���A�����j5���E�	?�/�;���f��X`Uj"ܭ;��i��5��8mW�ZE�	?��}e�X�}=��j{����F��_P^�A�qHPP5�%��v2�E��֢-�0U�B��J��+I��O�G�`�aw����m�iV�z��-�ғ>�>j�I�?7���x��6�4�^�=j"���L���I�Lk	?.�q������E��;;���V���O��7y�|��4d�_[��V��ŭ3�4�Ѩ4��J�ل�ZL�,�vF��a+���n�w�^XMU�y0��]"�	���,���s�cv��ρ/�����K��a$>�	r��7�}�x��=
nJO�&�����s�s�X�2|	g���]"�	!�/��.0�S{�n5���SrRf�5՘�&O�a0FBl&\�ϝ	��'XO����&��k(Me=u�&��k.c�Mn�Қ?���M'zȳw�f< �G��bM��K�?f�"c�S�YBk)�Ys�G��d>n�k��D�k��bcLq���'l�� $�p���&dD��:VR�(qYJ��5�2F�N�8��p�S�Co���=��yF�����5���$%i\Li�7����ҽ�<�� �ȣ��agP��"�Q���P����v��Y�,�,�05� ���,,�jv)�i3I=��n�X��(;n�������`�Li��1���������)�74�6~c+�$���}��}�\J�D[�q�E���ԟ�$�sݮ&�r������.���0p�X�G#	#���0�/����0ܱ/����0�s������0��`4�����{�\��?�@ $퐘�� ��7�̈�YGJ�Ue+)U�&��H�)�'��
}�m��r�T�.��iQw�|��$�;em�v��$��i[�+��K	���I�H5�s�O�)�&{�N��`G\��)�	�C�~Zl$�4���(;n����Z��0E������b����=wQ �����d!�Uj"܍�H����J�H�=�.w)������� �Hn�H�L�r�w�� b���t��)]Y��`!�5�'	�c�R���T�v��cD��a�.M�<M#y��'��v�LOG	�@I��fDJ���e*�����Ys$l����w�>�T6��aHw��yF��q��D<�-@�� 7���(;n�����:.M�<M#�{�f ��J��ݑm�wd[x��H��E��$��>Ei3I=�n�X��(;n�������F˓lM�>O�}clM#�>O�}cm��>O�}y�:0���X�a7Q&��-+݋�v�	����GȪ�E��F~>F�]�
4,�0PUj"ܜf�f�O��/{� )�yI"�K"�XI�ob��q�a�����Q���P��j��@�	|�?դ�"�gdjH|a${_�N=e���OT#�t�6G9�x�v�ن���f�����I�3T儮���0�����ij�
�sGhy��hGR(0�9ۗ&؛����7?4������Å��� X�I�H�n��0�i9 n~i�%�����WDVw]"����ݼ�a�g@����K�9�������0�~��Nc���R m�cD�Q�Y�8���v�LOG	�@I��fDJ���e*�����Ys$l����w�>�T6��aH?�TmVas���E�,$>�_`�+H?���H�"����5}�ԭ&i!�r�j���2���Pv��aq%3C�����ecc������Jf� ̈́�����	!��;em�v�Q�f�e3�5&�	#�,��.TmV{���4?����� W愬_��Pa$s���i��W@f{.:\r��	]1Y�`O�r�3��L�C�&��a0z�!8M���˘�M��F�cE= �	��C(�� ����`f��(�YJ���e*���\�%;��B:���O���rR��8����	 \dQ�R�H��R��2��a ��?�XH���5�_ÉR������n�X��(;n�������!�r�0���X��(;n�������3H2����X�a$Zs��.u��E�We��sl)�h�����h����� ���<�qq�G�"�Ú�Յ5��%��<�hx�3���|�3��g͡���ZL�,�vF���H�OCt��Ff���7K=V:_�� b����@%�RFa$s���CC�g��7�WDVwCC�g�I�E�՘�&.TmV~�p�	��'���a�	�1�)묡5�t���`���̦�f�7�cE?M~R[���He ���B`z8LL�2"Ue+)U�8��VP�˙#d�p�GS�|)�Z���C
A�u�k�
f�Q�DR5�aq��\�&�+H����5�H*l�J�|��/I��\@ѐ"��I�E����"S'��5�Ha��Jf3H�a'ᅦ�n��&�� �}A�E����2�E����s�zV���_��ayyc�ԟ�������|�������ԕi3Ij�O��3��� ͼ���Fȁ�E���X^^X�5%ZL�,�vF���I��k�!ф��_���
g2�e�NT�J���v�Q���/I��՝� ��>t���Z�]qY���HÂ9�j2k�4�K7 O�_��3I.��a0A���1�(qYsÄ����D�?<��4'��v�LOG	�@I��fDJ���e*�����Ys$l����w�>�T6��aH2����o)����^K	���o^ü�]����_d�`/�E&��(�Ɣ<�u���{Tf��o(ұI���
 ��䃬���	 \gc�����V�4�b�����2���Pv��aq%3��3ln�1���������)�74�$�8�V8�I�����$F"���m)�
RÛ�S��J��U��s)�i�ͱ�μ�}٭��\gc�����V�4�)���#0�9����q��~�~n���%��� � z��c�c�MG9fm��/���6��_�������WDVw �] j��D0�xF�8�He ���B`z8LL�2"Ue+)U�8��VP�˙#d�p�GS�|)�Z���C
KQ���5�wɮ݄�Ԡ�5�!��y���k�*��aq+H��0��*)Ջ*(۾��б���x��5,$q�������ZL�A�'��1���������)�6�0���2���Pv��aq%3�f�OÌec�����q�������U��s3H��������i?�K=Tfi��4�ۥ��3��WDVwY���H�$�v����g����Fۖ&�F�J聊�� K= X�Rf�16�&+	����&�	�h�����\ǰjo�`6)F��"��|y���P	;d&'��� $��3"%VQҲ�YC��Ue	���6Jw	��u;�E�|�0�нY��!E�'�`Ҹ~,
1q�V��;yIV�o��	�_�Z�����~��x��Jfz����������4��~��	{F&�:�Ef�HQa��+�����V�-��sz]C�Y�^���
��Ui1XI�D�d���7M���ް�8�ƕ��2�E���Fa�%�>��Ô�Xc�x��O�ǟI���n��C�u�F!_�:�/��1�Gm&��C��X���a7Q�󁊑����Q�
1q֓4�)��� C	��I0��8�H�{u�̀��!.�a#Spq������C�B]#����S�PP��j��{F�6	`�Sr���
w�^�`=����1Ƌ��	���P	;d&'��� $��3"%VQҲ�YC��Ue	���6Jw	��u;�E�|�0��qZW� �u�qe��	 \gc�����V�4�f%�ջ�ecc������Jf�"償����	{�C��I�Á�б���x��5,05�V�-�8�"�gdjEG;���{��Ķz��a+�+;�-Q���챝 L�cEq���b(R@ $퐘�� ��7�̈�YGJ�Ue+)U�&��H�)�'��
}�m�h]F���m�TE#]v-��}Ui7Q���SeV�弹�T��� E#V�4�D�L�B�a��Jf3H�a'ᅦ�n�߫d@(�_PiQm�=���n`"͟M�����������@�'�v�/�������Υ��ʴ�6}7���=,����w����ƻv�7����.u,NU�0g�������M�ZW~[���Ȟ5ۿ�xoդ� ��O��7�3o) 4Ѳ iQ}����=1��ZL�,�vF���I��C�	���3�h�'1����J���v�Q���7�gd@)��"� �b֮\Vj=j�0��r��/R�M�����Vb��	?M~R��4Lz�V\ǰ�$v#�#Dt6Q��k���[�oE!�N�	�@I��0	3xLȉU�t��VPⲕYBk.d����p!N���j��9)*6[�^۰cb}��}���4��d�%�+I�O8�V�:(����S'��cXI�q��qj�H`��Cմ� (�vZ��0���x�V8\��żD���jXpv*�na�iS;#RG:Y��� ���	]]��`���jX~xu/Yn�{nդ]1��+;�H���#�"�!�N�	�@I��0	3xLȉU�t��VPⲕYBk.d����p!N���j��9)?�f(�X��7��դ� �G��C������������Ԫ����Y����a7Qn/�4��z�\`(�w��(�nq�X.����/��]{��F9�ƨ	�R~K��k��r�i�/������ ��OÁ��^�G����^�jX4��z���n}fQ��%�)}C�a��\���N�%"͂�7��:���� ��(���g������S��-l�[�7.��c�@n����u���"�gdjH1���~i�4�3�iФSa$}j~��x����m܀:��s���m 8�M�� 2 �]�{Hq��#�B��'l�� $�p���&dD��:VR�(qYJ��5�2F�N�8��p�S�Co����>%��i��vEn,�۰����\�b���=#�5�>'l1{X���{��j�j%3/4��$�8�򺈣q}A�p<��nI�a'უ	#��8u�]��o���R��e��r�cZ�԰iV�Z7��,�|#Rf����H:�J6���A���9f���-��Gҍ���P{��Y�Ԫ��D�r��H�n�	{M���Z������c��o�5�/�4�c��r��A�$`�����!�����17�ZF� ��%&+�Z5�\/�`��T��\�u�b���Z���XI��Y�7Π���}���TJC�����7�h�j��20UZL�,�vF�\����Q�A�W�{c2�Y�|o�&�C�	��Cx�hޖ8���`��)��R�1���a��a_ZT�G�Ҵ��2]Y��`$Մ�L��	��&�Lȉ�YBk(Me+(Me+.c��c�3�B�j]��S��#�``(R@ $퐘�� ��7�̈�YGJ�Ue+)U�&��H�)�'��
}�m���������G��Á��v��@��S;�d{�8��`���Jg���|�R�Bs	�P���s�8֢Va�.�}�;KQ	�'� G�?sR�J��a>����������֢Vey�Qa'უ	#��8u��l�T[{�x�Q��C6� �$}(��p5�� `嚃���H:�J6���A���9f�R���ʆi#1�G�%�]6>�nUj$�LV7-��Q�0�,��ҭ��MʼZ�䑃��� �_S����ic|����/��k�_����&i,$�8�+��_�z��+���Q�ךM&~Q!�l����Z�ԁ����������I��	��|a6)�tBfDLz�YBk(�YBk(=���`"G�pg*�Ժ	�.�@]F���f/�E�E
C(�� ����`f��(�YJ���e*���\�%;��B:���O���rRHz��H.�t;�u����[�^�c ���8$^^�$��i�d@Ҥ.�t0:�i3I�={��ܱ���%3Hz�Do����_�[�^�c ��%3��\����+r�&�K��7�$p��Y#�FʭD[����O�#vax�����iX�߆��E�����_ZT]�8b���~Zl&�"�����l�x�	 ��Ƃ�E�����>�߮N��������lt~o"F2��i<g<[{�~�Rf�9����,a�n=��,a�֢s������a�'�V�7��N~a�4�$�&����PiR-͕]v�t���*�x��&iS;#RA�$�r���y���S�簒9�z�)����� ���DC�"�!�N�	�@I��0	3xLȉU�t��VPⲕYBk.d����p!N���j��9)�m ��yV�4��|E��`����t�L��O�a�j!9��@ �s�8֢V`$.�}�;KQ	�&�#Y�$�q�H`�OÁ��+��7�TS;����vjr�-D[�qX���P����7�
_��_x���i1XI�`��H��]cW{t�����԰}�j"ܼ��ּ�,TS6��5;ԙ�0cm��Gҍ���P{��Y�=�t�����o}����x���j5*��Q ܨf�3�|�^���c��V�A�t�cpr��u�r��*��tܫŨ�nI1}?��e�'�<M�V��7�,pII�b�F�+�����f�I����^9�m*Ӵ_Pi^�]� �nV�X֮���}���O��!�����%wQk��Q}A�x3Uj"���I��O����46����j�w�mӒ T��0z�1�Z�p�C��s��5���jDfP_vD<���ȩ!���V�4��YL�Hta7Qj�-T�(�]�D>8x�o� ��K]�|0W���Z�V��J��o�
��ZC	 ����&i4���a0|�&�`!�M��I��	���:!6�	��c�RWYBk(����P��YA�e	���e�{�|�NY��ȑ�ܳ�=���;c����E
C(�� ����`f��(�YJ���e*���\�%;��B:���O���rR�r
�/�H.����Wt�B��X�}�S=�q��&i ��=�z�D�`.i�I��0���7�$u�b�욙�ÌUV�-��4�L$��p5\=>��}�H]����jg�qD]��Hta'����i[���:ȇ���En,�۰�]���((��Ϥ\�kJ�����_�H���jX7�h��Ui3H����a7�)��z�� C��E}�(R@ $퐘�� ��7�̈�YGJ�Ue+)U�&��H�)�'��
}�m�v�d[v�`yV�4����n�݃��P{��j%2� =�;KQ+0�����̯4�+	?�<��(�_Pi[����<J�����Z��$�1���E��x8����$�0ta$r�� �����m��W�jX>�n^C5�-K���Z7��,�|#Rf����H:�J6���A���9f���-��Gҍ���P{��Y�Ԫ��D�r��H�n�	{M���Z������c��o�5�/�4�c��r��A�$`�����!�����17�ZF� ��%'���-���0r��I�G�	?:6�st�U�h��ҷ݁�u��E�[�Ɗb]�]��B)��UZL��$�/�j�sCi[����5p��߶��	*]wI�ŭz���}�.uF�ҭ<��Ch���ȇ�ҢJ� +�a�V�4�)���1XM�Z��U �+���a⡼X4oKH�a-]�|0W���Z�V��J��o�
�ҳ4i=l'�Ҵ��Y�Y��`$Մ�L�)	��	?�a0o�&�` �? N�ME���P��J�(Me	��5�t��5��\ǰ�pa�,vo�#���;q���.�����N7�l`F��'l�� $�p���&dD��:VR�(qYJ��5�2F�N�8��p�S�Co���2#py�8o�X�i�
��B�	�'��ZLn�PA��v<c "5��K	�#f����]�����J��V�4�i����60%3�ǜm��	��)���q�Do�)�ǀ��8ۢ7�).�S0�i-XI�Dn���E���w��$(��n����D[��a'�8ۢ7��ZC�o!}B@����E����$�'tF��f$Â蘪r*�nF�L$�'tF��B�	���&*����e��s�2�V�o�Po%���GѨ��ZE�	?�c�DX�X�b/�4����
�D[�e�^Ɇ�V�4�)���L�n���+]/���`A����KV��a&�8ۥ��侙�F(�`!ĺ�&�5:C	�m����J�ф�ZL�Bl%r_L�DjA��)�Ӷ��"F�-x$�W]�t��}��a8��S�1��E�&i ۫1XL n�hNDǬ��e�{��ؕ2F�c��60��7hBi�2�@I�!0	=&&o	�*������VR�(Mȇ�S�N#��>�-P��!�'�������c�� *�y�����.�*�y,�82x� @����a 7Da��@�����ZL��?7Do��	L���?7Do�&bD�F�)����
D�q�)��L~n�����;�L���Y����݃װk��6��3���#��Ũ�sG�
X��Ѭ
����4�&�1v�/��k	�x�Ht`�,Y=� ��x��1����x����K�O���?7���RդP`��%��i(��a-`a,�ZEX,�lty� �p��Hr�e��Ѓ[">*�K`���v�iX,��,�p��I��e�,�0�LA��q��-1]g��E������D���xbX!zg�VD)VS�YsR���.�ρ�-��b�������U��"�	?	����c-!�
��A_�*�߇�U��s��a'�1��#�3a�����r*�nF��~��7��M܂�"�aȨ*����E���(��U�Y�
d}����ZE�	?�c�DX�X�b/�4����
�D[�e�^Ɇ�V�4�)���l%uq����"ԇY���!�jX>���$0a${W���q��� ��H��	��R�F��=ܥ~�`�uyo�7��v�q��)��c ���.;����`?g�)l&c�t���laHea7^ d��xL�r�s��f�B9�dZD.ږ=>�s� jX`"�t��:O�H�a"�:0��I�Hp�_�`?g�#RBlt�+.���AT����a0���|��	��;�H:ȇ�& ��|!?�&=e!:�YN}e�{�Nge#����2ƉGc2�Y���B�υ!�N�	�@I��0	3xLȉU�t��VPⲕYBk.d����p!N���j��9)Ņ��-��>>G�J�o[�d��\@_PiY��A��ԙ�T����3��=J$��L�wb8�:���L�f�ea'��o`תȁ�[�.8�=����ni�i^i�$�84z�H<7a$r���J�o`v�����H�0;^-D[������dC�k�i\-���6v�l��ecnb-�TMo?�6�3u�c��4�Rg��,p4c���I�O�=ُ��֑f��<^L'�⾤4��,��`)�ԢA�!����h1iw���ƌ�2~C�7��!�>4�67@��3��g�"��3a��Rg�"͍�{���������]�\A K9��+���I�G��X7�[m�g]C�d�n�	���p;T��n��f�aʁ���ר��,��:G�ҸZ5�\|l���\�p�cZT���d7���&i�I�v#�#�n�K��w����E�Y��Vu��q&��Մ�9����?�� #��=�Y��`!�t���6&?<c  ~n Є��	�1�)	�P���.cߢs;)�vG���M�x� C���'l�� $�p���&dD��:VR�(qYJ��5�2F�N�8��p�S�Co���2�������T��PÑZLn�PA��v<c !�\}԰��0�i
m*+�7�;/+I�IYP�����B��H�̭dC��Je�P�%��Jff�f�O��(l`Ť>N�a�
��"�Q�ls	?��I�9R�xCEV�-̬ea'�C���n��ʖ��r*J��`��n]=��[|*�y,�2>�@�(l`� �a'����K����E��xS����U��rJ�8�Aa��h�i3H����s	]\`/3w�\����l`9B��E ل���)9VG9L�H��R�c횪�Hn�TM�����&{����`��H��g�&iS��I�7�������7 M�nP��? OeM�r��?��H�*L�f��uf+	��9I���&��YLz˘�����D@ә�He ���B`z8LL�2"Ue+)U�8��VP�˙#d�p�GS�|)�Z���C
G%�iQF"���Id@ҷR!O ����f��cOt_�L��H�a'�	!��;em�v�Q�9�YL�Hz�H1)�-w���z�=~s,����j��~��=�9�|���fz��I	����F���n�1�����3��0�9�c+�z��^�c�S�� к���B���v���L���� ����BK�'�DǬ�=e	�����=��;݃�5v��4S~��4����BK�!�N�	�@I��0	3xLȉU�t��VPⲕYBk.d����p!N���j��9)$>>�1	B��*���?t���䳰���N����3IjҢ�7+q��g�a��i 7�b/�p4��f�Ё�l`JfV� i�ĉL�z�b�L����&4�`3�).�S<�iXI�4͌�C�(�j�aȪ�E���0�� i�ę+ �(�j�aȪ�E�t:0�� i�Rb۹%
$��r*J��5c�|�nVNF\U�Y�
d}�L��ZC�	?l%���U������@��wu-j"܍�����Ѿ��uۮ�^Á���!�.(�Y4����U��a'������E��F"��J��)�_P���E�$��Aa��h�i3H������1��C������a$3c
O�$�q���Խ�2�D�Q<��=�/AEr�=,��N�a$9��$�C�{�K�s�ȴ�u�|u,0zUSrRr�%D�.�@ɸ�MN0MĤta3֓4��	��5$c��������:�K�%�9�d)n�)��w )��ww�M�I�@ә����"ʓ4��Y��`!Oq����l&4�b�DLz�c�P��<�.c�|C��x��S������ZC(�� ����`f��(�YJ���e*���\�%;��B:���O���rR.+J�|/�H�,�ZL�z�7���S+,��$�"7a/`ש�mw h��ⱖ�-�f���x��J丗�����f9�x����5&+1�XpA֋h���xѤi�{�o��� ��yl8 �E�O`Ѽ����`oI��s�u��+Ph�4in��y��=�H?�A�h���7�v�,�1Y�3a��B�'�h�4in��y����ُË���O`Ѽ����`oI��u_�-����F����W�!����1�qP���7�v�,�3Hw���yE�agPi[������92�&iS;#Rr�$�r�������5UN�V�TM��0��oP2n0������q�G�mH�a3q)%l%Dڐc���~�g�U���:����Y�`n�$�Hq.�!���3H3����AЛ	����sq?!?�&=e+(Me!
˘�&5�>���D�F�C ��.n'�!�N�	�@I��0	3xLȉU�t��VPⲕYBk.d����p!N���j��9)���y�8o�X�i�h�PÑZM-.�*�y,�82x�s{���tF�'������yga�����yo�#�l`Jgz!�����H����!�����"S#�0��7���!Ipw��sH�a'��&�z���r �����nk4�V2#v�:���aԜ�a�x�����Nf0�ny�h��9���u��-����cl8�����Ot��b�/��o<m�&i,$�7���60b� ��U9Z��8�I�o�#�3a����U9Z��/%�	?�Do�)0���B�aȨ*vZ��#�1���T�g`)��j760V�~�OÃ��ۨ���E��xS����U��rN��y0�
�f�e3�5"鄮�0����ZC+	60����E$&�D7�s��)9VG9L�H��R�c횪�Hn�TM�����&{����`��H��g�&iS��,$�r��X׽l3<�yg`�����H�*L�n����AЛ	��7��	�1�(qYBk(=���a�c]����������ZC(�� ����`f��(�YJ���e*���\�%;��B:���O���rR(\V�b/�7�D������o�V�4�D{%2q�C�	?�]�R��U�%�1���>c��J�T��Z�V��{l�+�����i3H����0�Џt��q�Y��` ��	�	��#߀l`{��"c�P{YBk)V\Ǽ�^v��C�T�F�G� ��.�'�!�N�	�@I��0	3xLȉU�t��VPⲕYBk.d����p!N���j��9)�{���p� �����T0�V�KK�
��K;���]�����3Hy���1���b�%;�yZL�,��l`Je��w���)����b�L���c �tF���%��Jf�!�	?��1i��8PÑU��r��O��s1&xa�G �r*�nVO�~{��n���T0�T�]v�aj"����-�A��v�F�w�ci$�"7f=�E��߷Ob�%;�.�͌ G���sC+���`Ҽ(,7��	�U�R9CJ��X7�̡����7��~[����H��OÃ�������E��xS����U��rK��p���L4B���YL�I��M� G����
HLk�(�&�R<�M�͌)L��!G9LLl`Sr ��$a8��;[�\`#�$�n�&5�'z��%����Lk�N�]�`15�v�ciL$C:GF=i3I	��1�<��������>���G8A����AT���]Y��`%��b�p�&=e��1�=�`�yF���'m��v�LOG	�@I��fDJ���e*�����Ys$l����w�>�T6��aI���=�Lr�aqvv�/�5Ha�Ƥ�"�	? ���h�o�э�M� �C��ZE~>AT�Ѿ�e�J��l`z4�l[��������!�x3c������la�ZG�	?�I
��a��%�}��F6�60T0�i-X�q��N7�l`���M�x�1��&��H��_���{��#����㤈�,6�HP�&�F�}��m*l`���IR2W�cUT����V�4�B��V'�60	ƄضL~x�1�	���&dDǬ�ڲ�k(6���e+.c�1w�yIGj4�wj�xl`���Ix�
��ή`�nS�60	�HO艏YH^����j˘�M7۵�;3Li��1�	��!��l`�l&�� �p����*�YCe	�����=�W}��;PQC백�cDA�m�Fνv�Z����@ $퐘�� ��7�̈�YGJ�Ue+)U�&��H�)�'��
}�m�q���A�E�_P�W�G��h��7��c�� �@��>��U�8h��h�o�я��(��}�F��xɘ��C���x9���sy���'�&=��b_դ�"���V'�60	Ƅ�L����c�b�@��>�Lȉ�YA�e	��ڲ�k)	�\ǰb�����^әݫ1�$ܧ�l`r��	��~��Li�l&o� ����j�YG�e	�����=�s�T�=�����x#߀l`=�p�&=eu�1�M��<����M��A��2�@I�!0	=&&o	�*������VR�(Mȇ�S�N#��>�-P��!�'+ym*.o�ah���$85�8;`��By%3!������zBS0�4�6~��lQ�	��c�@i���r��
�8qZ��+%~��9�w��s� j㙩j"��Ό����f�e����4;��s�*C�0�".%��e�8|p<�T��Egt�6ash�j��^Ҹ+�_�>uiXI�Mqx���?]�ȁ��f���r�tf�n�
�$~T��Eg`!��~3�((�N��Z�爻V�4��$�5_���i�s����~���ԟF-��*�c�lV�4�Vb��	3W�!0�	��Bl&S��̈�����P��8VP��k.c�5?wfPC��t3OAv���!�"�!�N�	�@I��0	3xLȉU�t��VPⲕYBk.d����p!N���j��9)dl<(-�B�j�n��G݁����HT��'���{�,�e���ZL�}r{�S5$Jd��Lk	?
l��|M�j�����5r�E�Z�,p��ⴑ�I�`bL$�^X��5w�X>���nq�Ht`��Y#�F�����=��,���A�H�Q����jw�@��5�UU��*�Y�\#��.�p7*5
��q�@\��S��/�<J����/��zE��2m��~R��.Ԟ�)��r�������XZ�nW���+��c��o�5�/�4�c��r��@\��b����!�����17�ZF� ��%#��xZ5�\/�`��V�4��~<Ew�Y��s㻜����l��dA 5Nf�C��*�$�/�6>� �r6Uga 
�&��"��k��������$�5�pj,p\�%J�f����V&s	��	3W�!0�	��|a3"&=e+(Me=u�&����1�8Klw�i���r���)�tBl@A7BDLz�k(6���e�{�OAw��;���� ��b~R@ $퐘�� ��7�̈�YGJ�Ue+)U�&��H�)�'��
}�m�!��m;Z��M/�Pj㻆����pk�]�}�;W���2Z�.�i7�����R�v�4��Y7�!����&i
d?���R��Jg�.၉���;���;�D�G���a'� ޱЎ^X����8h�7��vD<Z��.��
ҷ�5,v*��7���#���v�2��� ��*�8|�v�]�,_,�� �ðܦ
դ�a'၉0�9yc�WY�����5׀�1e��s�t`��W�0;J��B����|���JLV�`39�_�W^�&ю@�q�r��A�ߒ���)��|�ᅅ���H�a'����{����E�	 ���CK�pw-D[�FVga���TW�wʚ�iڲ*A��ZT]�͕Y4�
�I�LV~?����}�9Iɨ4��ˇT7��@MI�b�݁�͑+I�E���Ԑ!����n0����I�w	�ҕ$.�B9���*HM��J�1�IU����	!�/�S�:@w��DA���'l�� $�p���&dD��:VR�(qYJ��5�2F�N�8��p�S�Co���W=iQs|a�X���G���8^�/�7Ɠ��!���7�Q���5*���JF��Y�c@Q���5*���JF���0ƀ�'��&jUUIL����j�FO��LԪ���)��{�������UU%2R�#����&�^�U�X�o1}C���no�'`��t���Q�l0e�(Ң���\�_�.� �q�� ����_�ž4|]�� ��h�ҭ��\e�a'aǧ�4�6\E��Y
5$�3/��Y0���i����7�+��R?�y���1���ˈxJ�4y��cY+���&�/?uU�%dE����/?|M�S%bF��&+	?�Xk���o�)|�}�8
_����v��3�{h����	)!�H4J��~���f�����J���r��\�^���I�ZA��T�"�	?���8�7�@ �6Ud@ё�� �H0b۝X���{|A�l�ȃ��!M�Zyj�"�V�4�)���l&~�6�0{X�)l&@q�%�ջC�"����S�R]�^�_P�)�JL�)n��a0�XW��Bp�&=e �˘�������#E3W�rD��2�@I�!0	=&&o	�*������VR�(Mȇ�S�N#��>�-P��!�#�P�$A}���r�b������A�H�Q���ے*8m��a 
�&��l:N�x:�R�v���"���)��� �$}(��v����x���j%2�3c���t�����o}��P{��Y�Ԫ��DyeJ����jt�����m���{��Q)���~�[�d��n������ `嚍J���CJY�~�����K�7M���G4c�����nV�0��d@Ҽ%iI�a1m�E��D��Y#�FʭD[�E�	?����Ӵ]�\]�}A�D�<F����e��s��'��{�u��Ơk�{��)�o��5*��Q FWY�Y�����DS����TM�u�`|j��+Q FN#3�.E:˝e����"�#�a7Qk�u��D�8�"�	?�@��d��6��0�,��ҷ�G�Q�V��7Mʼ	�_ C/�?��boz��1�c�JE���X���_�i3Hta'�A�TJ�l,p
�$~Tx�6ﰾ��E�M �ŷ>1q�F�<�O ��7'�x����-h�(ߺ��l����4cj�v��b����TLH��"����&�ka�_|m������o�pi����t�Z՟:��5�N����m���M�U 5Q�v�&iS;#R�J�&��ᄐj{�34�3O�H�nK��f�X��&i�Vb��	7$&�`$ư�	��.��	���:!?�Lz�-��5�8��5�VP��k.c�`�m� eGn���kݨ.S�]�ُ'�i	��G,+��!?�&=e %e	��Ys�P�;7r$ �'�� j"�!�N�	�@I��0	3xLȉU�t��VPⲕYBk.d����p!N���j��9)>����l���۰����,pu�݀�w�h�5��f��|}�|MJ��)�W4��I�>,&�"���	"7�V�-��4�6~Zm��#��@ղ���]�$q��!���U�����F�楄O
�I�i��$~���݃J��7�}�J��*��^�eb��\��D�]��4c�%�W\m15V�4�)����$�T����XL�����)
l$�r���?��
n@��q��G�	 k!�'=���S{�ã��$7�s��4�+�1XL�t&�`$�^ ��DLz�VP��z�.c�p���>)�����Ɗv����q���'l�� $�p���&dD��:VR�(qYJ��5�2F�N�8��p�S�Co������4�*)�_�5s���H�]���]�f��E��o�}�zΝ����V�4���M�o��p!��)�C�"�p�翜j�Jf�!償���WQn/�4���Q���OÁI�ҷ��G�S�,p`�KQ���a:�;��|I`+��E�^��h�����E��ҭ/YӴ]�\^ڙ�Q6vդ�"�gdjN{	 �!��a�l�o��E�	#�;i�C_� E��������˫1XL����NDǬ����=�S�v���D�_� ��P	;d&'��� $��3"%VQҲ�YC��Ue	���6Jw	��u;�E�|�0�={��v*ר��$@(��a [�d��+I�HC�f��5�A�H�Q������>f�I������t�����eB�W}�K�R��ĠjX�V�-ˡ��%��u�2m��~PNJC�u��c��V>����׃r�դQa'����H`��tۡ 5�԰�Uj"���Hw���!}A�E?Y���[N��W�v�e�����yPF��Ŷ�Y#�F�1G�����*�=��n���[���ŭ���k��i3I�Vb��	5����4Lz�z�.c�5?���#DB�#�B��'l�� $�p���&dD��:VR�(qYJ��5�2F�N�8��p�S�Co���=iQr)�\�_|��դ�$!w�ʚ�;a.=%33I��O��$�*�6ǋt$���,[J�u���-���$�/�a�+I�E��1XL����M��I�O E�'�DǬ�����P{Ys����2�S��R��Es�)�v�LOG	�@I��fDJ���e*�����Ys$l����w�>�T6��aI��PP[��l}�(�)5,p�0:v�� ��dA `����\��)�Z�t	L�f�a'�ф���V�-���(����m� �ð��`�"�l��*�G<E�5�i��4��!�xq�:0��{�.�>��	q�)�{t� ��*��Y�"͋l���5��U� �^����ܾ�s���B�vtR@V-}��fYAq��դ�"�gdjC+	��aga 	+H�a+�-������@>V�E���S�۽e��V�����@�}{t�G;	R��L$�r����z��.qq�����x��� �v�i3HVb��	<�HNDǬ����L�k���)ƈB��~�?)�v�LOG	�@I��fDJ���e*�����Ys$l����w�>�T6��aI�1���u!�a��X�0]��bߣ����
b� �e��o�(;n�n۰�^�!v�W�"}Ui3H�N� �$}(��w�P{��Y�=��H:�J6�����x���j5*���c9/�n�u�>�m���=��,��[�d��{��jw�@��5�URS1�Hta'�|�n�(�_Pi^���(��Rý��b���E�t�g���[b�sP���%�)}A�P5,g4�6q~K����d�1�.5B�����,����)��|�ᅅ���I��O��0r�pA�J�k�_PiV�ۦ�^���Q�V�g|	�O{դa���`W���f�e3�5"�	��Uj�Ez�b-+r����:0�=Cx�hޖ8���`��)��R�1���a��a_ZT�G�Ҵ��7����I�!6&j�&�"c�Qme	�����=�v����݀�������߀"�!�N�	�@I��0	3xLȉU�t��VPⲕYBk.d����p!N���j��9)K���m�Zv��:�z����1=7��[�d��K�-��Gҍ�IL��i$�-��Gҍ������Gҍ�XN��X5w��U����Z��E�Y!�VY�YL�IL���	q���`{I�a$s��v���`Sr���$&�q=7��Ho�>���I�7���:0)�C�ސ��������P	;d&'��� $��3"%VQҲ�YC��Ue	���6Jw	��u;�E�|�0��#i��\��B�e�]g�դ� ���Z<�S/(@ ]�x����ܵ���=����9|ƥ���|�IL�%3�T��VDj%�)�L�b�������WuF���J�k�w*��P���p�"�E�tY{�R��ĠjX�B���׸ɴc��f���������x+��xaak��_��~na/q ����J�h�p�1����E�?XI�`��72WuK���^�W�?��e�'�<Z��.�F_{դa���`W�9դ� ��O���5x�M��	��8.S԰����$�2�n�`W�9j�f�e3�5 ����s ��N{1,���S i!��{�	�U#Ʉ�����VA�Gc3�t��6������/RB%Gc3�t���<Y�8�MrP���IXJ��g��տ��i�$�r��g����x�_Gc3�t���I�CM՘�&M�	��	3W�!0�	���:!3"&=e�P��z�(Me��1�0C��_'���������DD�Ř�He ���B`z8LL�2"Ue+)U�8��VP�˙#d�p�GS�|)�Z���C
E�$��vu�J�k�+�@l}dA \֛*,u$&�_E�4��$�&�LZ��/����[/ ��t�����eV�-̮9�����Oa�z�}v"�x�[�d��*�nI0����[�a��W����(.Ml�x��}�A�H�Q��Q�h������%oa��a�����}J�[",7�n�u�>�l��E�Z��O��S Dn �<��4[Dn�<�V�-��A����VJ��� �$}(�`_a���A�H�Q��Q�ni��a0�g��!DIp�PnHLȉ�YJ�����²�*�-���Lhz즪:;�4�3O���q�Bll����Lȉ�YI]e+(���me=u�1�K���v�QO���f<��	��!O��a�	�2"c�QҲ��P{YCe+.c�]
�����r8�'p���KXNDǬ�5�1�CBv����!Q)�v�LOG	�@I��fDJ���e*�����Ys$l����w�>�T6��aH��$]��waw)�a _v�i3I���SP
7{���55�2���OÁ���Qn/�4��4�`!���nIQa'�!��n���X�o{K	I;�5,TM�Q�e`�UM�$&� ��E��iZLV�)���F�}���F6���(�Բ��޽��<`��PۦSQ�a�V�4��~]A����!^-?��^sJ�� ��"^�~�h�b�G���U��"	 �S	U ��n����_ ���U����!���h�� �S	R��,$�7���^T��k��p�C��s��5
�(1n�h�x���VDzդ�"�gdjLVu�"�H2����}�x�o��R,�KWs_�>!�A��"Ҥ>[�¾���O[	���&in��a0�f$&�`$�HM��A7BfDLz�<�(Me%u�&���1� �����X�S���<�#DB�"�!�N�	�@I��0	3xLȉU�t��VPⲕYBk.d����p!N���j��9)47�I}v�]�jXH2��e�\^�i3I��Hw��g���<?��]f��O�C����<t���^Z�L�{�"�`W��j"���NÁ��}i[���X�&5����ŕ�E_ZV���x-�j�nec+#�Hx�+���!�o��+��ZL�,�vF�%t�����i��(:ȵ�!�4�L�,$LC��XI����)��=�	���q����!����n09�`=�1�Ww�zE�%d��>��������^7��a$=V��$����w���� F�Y� ;mz�.����e�\X��#���Я�A�E��5i:I
�M�<��7�s���LvG����"�՘�&MXM��A ONa0�XW��BfDLz�YBk(=��5��k.c��c�0���-RvG�� �E
C(�� ����`f��(�YJ���e*���\�%;��B:���O���rR/��I}v�]�
�ҷ-WR�漅�
�I�HL��-��Ly�ư�����n�(�_PiV��`ѧw)ga��U��r��"�gdjH�%t��o;v*�D;� �gadA w�HSa$��c	��@!ެ̪t��_�Y��`$Մ�L��a0C&�`!���������&���Qme	���e	��Ys�D;��I���Ƌ���A���Q6UUHqP�2�@I�!0	=&&o	�*������VR�(Mȇ�S�N#��>�-P��!�!�B;	�����E�U ]�l��|�V�z���};v:�i3Iʨ���������MD�L��	���5-D'0���BS$��Dؔ�B�'��Ե��}8����l6�@G5��/�I��%��EۦB�kt�k�a'a��Z��+%Y����8~��ֿ�I�E���ԃfa�8��A���S��}B�p�P��_P�Y���,7���J��]z�p����H�K����%�,�L�JC�G9N����M@W�}@^]g`
n@�ޓ4��Vb��	?�a0oJ��7�a0E�UTC8Lȉ�YBk(Me=u�&����1�H���G���y����
�b(R@ $퐘�� ��7�̈�YGJ�Ue+)U�&��H�)�'��
}�m��A��0W����	o���`W�9j�f��}�q�l|N�i ���l/�퀖�騔̼�~�bȃ_ t�k`�q� ςUZ��.�$�&���|�C�����n]�$�4���k���!��� �UUH�	R�Q�a'�'=�H5���?ķ�D[���I�	��"|�}�UZ��.�~Z�Ѓ_ ah�p�0�/�UZ��$���O�K�DX^Uga�Ĥ�E�/xk���iV����^��f�e3�5$�H�)�d���l9U:GF=i3H2�Y��`!�M��I�0�	��CUTA���ϸM��K�����1�(����QҲ��R��5�V\ǰ�9gp�B;��������+��1� �(M�` ��6,� �HM��%�'���YBk(����YVQme��&��=�����4���RN���4'`%���#�B��'l�� $�p���&dD��:VR�(qYJ��5�2F�N�8��p�S�Co����[d��l��9w� ��8/�πX���j�f�tG�k��;`�llzN�����y�c�S*\�XI�O݋"-�@#�``��n\�$�M��"�$`�*�nh��O�oKD[d�C��.Uj"ܸ*�O�o�	"�$*�D[�O�$��ő� _v�V�-ˆiS;#R�M����I[	Q6��t��aa�B]'C4�a�8�8��.4��M�L&n%$�H�)��ɪ��,7��&-՘�&�00��LQ6UUf�Bl&M�UUf�Bl&M��Lt&���YE��&��*�YO]e	���e	���e�{�w)�����=.�#�;��$N�T�cE7�UU!�B��'l�� $�p���&dD��:VR�(qYJ��5�2F�N�8��p�S�Co���A�$����}���}C�ڴ�������k���W�����v�;E�����a>��������{�c��A�Ԫ���L��H��O�A����l|�fN��E��j�D[�Z�	?�����a7Q�+5�B���["��v��* Ư�nN�.�$�,��v�;E�.�wm+q����PU�~����r��cZW�\�&iS;#RB�$���pq���6	qԐ��s�7��a$=V�}IM����԰XP��hR@F:ΰޓ���XoI�A�՘�&(�*��q!6'��l&����g	�1�(���5�&���S��=���;�G�k��y��S�ƊjIUU��E
C(�� ����`f��(�YJ���e*���\�%;��B:���O���rRH<�X_���!ZL�c���;���R��sJ���*Jg&;���;�MD�G��:0�����n�,,p
w
1�T]�N���J�Z��'~Ǭ&�"��� �p�m�J�Da�*�nN3I��O�K�5p^.%֡�Ĥ�@�$c�c�S�Q�W��/�pV�E�D����95�l�[y�HR[�Ri1kt@�W�8md�P�n�*���il[uZVB`-�+�W�r�PX���VD�R�.p�A��~��o����t��:)5�ݰjXMIRC-�Dv�&iS;#RB�$���pq���6ӚH]��),E �"�I��Hz�7�ta3֓4��'H<�F���$�u����d��$E�&i=�Vb��	5a6�v�a0��UU����Lt'���YBk(Me=u�&����YG
˘�!���A����}�挑;���� ��P�2�@I�!0	=&&o	�*������VR�(Mȇ�S�N#��>�-P��!�!��Υ���߃�ZL�z�:��S+,�~�&�"��� �}A�E;�,rp�UZ��$�ea'�l�����/ϛ���*��UV}�n�/�C��'����b�5,.�W�AoX�20UZA����Wga{B�fN�@Ӳ iSc "��*V�4��	3��e%u�:tA�w�G՘�&(�*��q!6&��l8��CUTA���ϸLȉ�YE�e	���e+)	�\ǰ7�B�;�Ȇ���c�Cc ����q�UY�\&�`%���l&	��DǬ��e+(���5�VP��8V\ǰ�i����w���cA"v;�F�H`���4UR;B��'l�� $�p���&dD��:VR�(qYJ��5�2F�N�8��p�S�Co�����{	���eW��7���I�Ha�0VX4	LÈ5���v,K5-D'0���zC �O@A�Jf簟|Ń�Q�UUZ�N`*�y�Jd�a>���KQ	�0���������?�w��o��Gxz&�S*�Մ���+-��(��;�����
$�e�����s�Ţ8��=mu����X���Z���E���XI�`v,Ka$r�� ����q �c�WYǡUj"��pk�v,�D[�Nb�ň��-�'�a'ᇢ�Y���+������52���V�-ϯ4�)���!�������?�zO�	����	`m���� Ф�t#��m��H�a3���B9�f��}Ce:A�	#]!�&i7Vb��l`���IBl&*��:�M��K����̈�����P��,�(Me՗1���ٕJ��������_F���UU����UR�O�C(�� ����`f��(�YJ���e*���\�%;��B:���O���rR-GI��5,��R[��]�U�Q}BH�c�����V�4����
�B���X�h�L�L�� +�W�ܱ����f�h0���턽���D*�c�o�g
�D[����OÃ�c��bװie�#�`X���o�]A�Z��0*�nVGF\Q���_�ҭV�J����Hte�W��r�A�E��|5����Xe�<���/��`\J�f��O����А.w4b԰�}Ŷ���Dg��!ⴙ�YL�IIM���	a�l��F:��B��/�7���1�IU��&z�f�a3��r��z� ل�����N��\`#������H6a",�3Hd����Cc ����L�>o�O艏YO]e	��ڲ�=�Pj�˹W`���Es��P	;d&'��� $��3"%VQҲ�YC��Ue	���6Jw	��u;�E�|�0���x��i[���X���઴������k�;���p��MD�a�b������ba7Q�b� i[����kÍj"���l#��o� ɪ]B"�S�Q�������HiaqI5�xX���(����fŕ�E����xg�q��]$﷎��Z��'
V *A�c�E݅ĭ&i$�.c��.5���[U������xR?X�U�4�-�jX5wHU���A}��1h���i3H����3	]=���N݃J�Q�H2��YH������B&�55�cA5�h;ՙ�N�4�"��V&s	�h���8���a�[c���#E~y�)�v�LOG	�@I��fDJ���e*�����Ys$l����w�>�T6��aH0���
1���*���4�^����Rc�}��}�\J�f��~y�-�)�B!��S0" ���X�jZ�Y�܇��S0�> {�v,��J���J�{���d�}p��b#Q�j%f��Ny)�^i=�$�0��ZC�K4v>�۾�.%V�-�����
2�pG/,p
�jX���Uj"ܘ͘���.����b���v�����rc� � ��(;n�����ư����X��H��]c}�F2� ���B��E����-��X=Z��0�Ÿ�-D[�O4�,$�.�*�����s�_P��{��c�JC�-����0/�/�P�F��'C�}��}�\^�l}��}�\F�UUj"����?���E��71n� `2�
�p?�D[�����cȆ��8h�?�7-D��֠Ά�x[uil��2�p�0�9y}A�E��2�2#-D��9�����w�{�����c�ƭ&iS;#RFa$}jdy���i�
���vx�k�����^�R@V~y������4���b���O�c��S!�Y����/]���
�t���#��F7�K3<ȭ�w�N�j�D��&i C�����c��S:���5�5,7�7�:�� �ܡz��HP?�S�r3�r�ޗ�^$(�/c�̱҅��]�����UN�4�6:��I���s���vxx�a��U:F<��)����=��I�C	#Q9����n��a0H`���4UY�	�h�����.cߢ.�(���*"�!�N�	�@I��0	3xLȉU�t��VPⲕYBk.d����p!N���j��9)
wr5^j�f�_���~�5���I�a'��J�H�2��w���w��Ҹ*��E�t�&+	?.���Jv X೰��x*�l�|M|�O�����	Q�JJl��puJ�f�e3�5"����Sސ�!�H�V<�IEUUN���o��9���I�?NC�`x��S��$0����Aa8M���\ǰW`�����HE
C(�� ����`f��(�YJ���e*���\�%;��B:���O���rR@G��
�I�C�
D�I�!ф���nRӽ�i�7���adA��n�=ԙ�q�l�o ��'b�	1����&Ŕ����nR2"-��ڲ�k(6��ʲ�j˛�8B����Qܷ"v�ŰcO�60	�8M��A�c �a���60�3""��<�(Meu�8������W|��nw,h!��iS;#RB�$���pq���6	g4���s�7����H`��#��@B�W)`'n@G�]�I��Hz�7��'+uf+ $���L�	�U�p��5�[Ys1�Dpg���=����E
C(�� ����`f��(�YJ���e*���\�%;��B:���O���rR.W%��aq����������԰iQtK\�&i%b	L��!N��V'�&�` �(O艏YG
�YBk.c�M��#�v����oz��<�Q$'�!�N�	�@I��0	3xLȉU�t��VPⲕYBk.d����p!N���j��9)��F���Q%�R>�l�^��J6GHgdC�/�5\=i3Hq��60%2J��T�H���i�$�E�auî�j�;n�Q�]����^"�c=��A�Ui3I�uf+	������j;>�g���1�)+.c�U=n�T��������E
C(�� ����`f��(�YJ���e*���\�%;��B:���O���rR��{	��Y�`_Po�'`(�������l�0u��f����*Jd�J���*Jg4�)��fJd��/�I��%��EۦB�kt�k�a'a��Z��+%Y����8~��ֿ�I�G�~
&ʪ�#t$���,r7Ѳ ��1kU�+I�M�Vb���l���Ą�L�Ҫ��������YVP��z�.c�
�㿢��`��� �7Z�2�@I�!0	=&&o	�*������VR�(Mȇ�S�N#��>�-P��!�!Ѓ �#����H��x(�[�� �'ǀX��n�����-��آMl..����Pk�@k������ �����kթ`��'=�͑L���@^����.%i3Hz;n�
5j�YeI����S2�Ij�O����6�%�C�*-�A���j"��y�9c������U����2�e
6��-i71���E�.K��x��[����CoS8Q��Y�#=l. �dFe�n�������A
"��fP�ݖ�L��t��迶[�~�,�HQ�F{Rnc�����4�e
,3�[��4��~;po(;n�
5�$�wd@Ң�ڎx�IŸb��vu����@�������ԙ�t_�em�v���Pv��aq�o =�(�z��r�_�-�#��h1���6 �x���� <O� �<O��<@�� <OƑ��M�c�3`�w�N�	0���H�c��1��0��	�a;�$`�F�6:���}�0a;�'y��N�#���c����F$`�F'y��Rf��O�� ���f�{u��x��ش\bȀ��������^�#=��0��_�em�vau�A���jX
v8���\rR)X�� ����+H2�����*(�kt�k�jX�c�b_� d�Ô�\�i�8%���J�۷��U]��h� �(�^,Ѭ=vw�"͋L�(3x(�[���"Ӵ�m�9_¿o��,5�qiضPqk�{�[e63�e��o�� x1ƈ��vސ�'l�� $�p���&dD��:VR�(qYJ��5�2F�N�8��p�S�Co���ZQ�ۧh��/�����4��;"	oJ��C�/.,w�Ѿ�g���#��%��q��$A�r�y7�}�l9ZL��Y��`$ޕUVoT&�` ��������YE��1��K�*�
�.1Ɗ�s��P	;d&'��� $��3"%VQҲ�YC��Ue	���6Jw	��u;�E�|�0��҈$	�*��W��k��oXt���R�S�ҷ�8_R?l�a�kaq*Q �����m�k.>.ԇ��԰i[��yk�XU��#���V&3��L�Ҫ����L���'o�6&��1�(����S�YBk(�YBk(Me�{�� �G�ْZz��9y���c~a��xx5������8��=e�{�w�۰$yF�x�'m��v�LOG	�@I��fDJ���e*�����Ys$l����w�>�T6��aIo�7a��5&iXI�=��ǉ}B@�<���i,$��^]q�Ȃ@�Ҫ���q˕�;�I�z�3,r�a�`PY�����3<Ȃ@��UU���i#0�� �o�ך�;"	 �Qc���*V�4�;�1XL����M��I�*��ިM��I��!6/ϛ��DǬ�����S�YBk)�YBk(6���`��ݙWH��Tҋ�c�ʆ+�G��"8E
C(�� ����`f��(�YJ���e*���\�%;��B:���O���rRb�J�n��^� �6���qD+߁w+��̾������&���W}���,05���4Z��,"x((���:Y��!E�'�`Ҹ>EBcHP5��������^�+��V�4���<��)MD�a<��$�0|�Vs֕k��"#��/�5�4�
�h��UV�-���,�vF���$��<�'4���Vb��	1�'	�c�P��=��� ��#��B��'l�� $�p���&dD��:VR�(qYJ��5�2F�N�8��p�S�Co���w=i[���#´���{��1D�a�i�$�xa/`�.��e�j_x)x+1<Z��2���N���	���$�VD*�c�o�B;���CK�#��]��ÃY��xٲ�+q󅔊��*.o�ab���YL�I	��=���&��0��ܥ~���`�uy�h�+I�a$���3���n�5��љ��.�\�jC��Y5����AZL��Vb��	2��5�&�`!
�HM��I�_c�	�1�)�YBk(�5���\ǰ���a�z.�=����1ƈa�_��ZC(�� ����`f��(�YJ���e*���\�%;��B:���O���rR8�+J���"#��/�]�8"o���&i �����ecc������Jf�F���-?�`.i1�$�8�V8�K�5�n�]��\����e��s3I�aLOv���a�R0���	�x�)SX��.�ׂ��J�ubo���9�qw��"�qRt���Y��^"o��Ɂ���aL�58�M�n�h�k�3I��O�M�1����A�w݅Ĩ=K�3/�RC={��;m��-��aM��Mp�� 7Q-���V�%�
m+we��ƚ8�i3H����M���S�lII�S����5?���I�7�&�8��fx$��{)�R�r���N�G9L������=K���� ��cD�_��^��x���P	;d&'��� $��3"%VQҲ�YC��Ue	���6Jw	��u;�E�|�0�;߫��H�H��-��$%i&˝�7�� ,�Y
��}E�	��ZL�B������ecc�����R�%3����x���ecc�����R�%3��ư���X��(;n�����$���}��}�\J��E��j"���>��x�{e�԰� TX�~*��ZC�>�v[�(x�]����"�gdjLvG�}��&B�8����q��$8a/� q���x����$�q��
k���!@Y�)�B���U!�7 >����D��!B�t�1����0����ZC(�� ����`f��(�YJ���e*���\�%;��B:���O���rRhU�R��J��(�/�H4l�.k��u���"���&��w�_�V/�G��c�I��O������n|�em�i\��-�ѕ�1QP��:�v�H�{�4)5��L�դ=a'၊�n��GR��V�-�8����?�����԰(,��8*�na�iS;#R�L� q���DS�Pa$s���W��4�17�[���1O�&i�Vb��	2� ��M��I��&�`$ܮ2"c�Q�YBk(�YBk(Me�{'�wоA�vdXC�v��Ɗz~Γ��P	;d&'��� $��3"%VQҲ�YC��Ue	���6Jw	��u;�E�|�0�r.K�ݰ�A�/R��QO�c��\h�N�j�f����-?�a�y��)n���Jf3Hz�O�M��ƚ;em�v�Q�f�e3�5$>0��Ԥ0S�~��EN�a$s���R�'�G:z{���R�� )���N��	#�!�v���R��0�0���_���S���#E2��s��P	;d&'��� $��3"%VQҲ�YC��Ue	���6Jw	��u;�E�|�0���lѥ���1�8��)c�qF���Dz��!ⴙ�)̮�-?"7�Jg��׻Oȍ���)������	!�4v>�۾�.%V�-��a'��0���}B���?�>���sK6s�1�� Q�,pa�(Ҵ��+I�E���ԅ6!H`�@��a$s�Wt�/;�DVw �a���a$s���Ga+�+;�5�&i!�՘�&M��8M���\ǰ��1ƈ����He ���B`z8LL�2"Ue+)U�8��VP�˙#d�p�GS�|)�Z���C
E�Ң�E��YH4K*(�_P<�[��aޥ��$t�����ei3I�d�ai�%3G�-��Y#�F��L��Hz�O�M��ƚ;em�v�Q�h0���>cȆD\M4m��Gҍ�Z��.��YL�HSa2��
d�N�0�9�-���f�]Y��`$��NDǬ�5�1�C˰N�ƊgS���q���'l�� $�p���&dD��:VR�(qYJ��5�2F�N�8��p�S�Co������r�R+���4�� w��"+I�HBgSv��S0�z��ZGB��-?�a�4��$�0��Ii���Pv��aq*�n`&iS;#RC�	��0Sa3]0�:G�G9LȦ����S2)�t@�gq��&k�d�q��9�fE0<�Φ�
_��
fE6� b���I��I����H�)���wHR��S2)����� 20������2ƈ�+ ſ؊�P	;d&'��� $��3"%VQҲ�YC��Ue	���6Jw	��u;�E�|�0��u�S6��/�H4wH��i1n�C��T;l>v�/�H4[4c���Q�D<V�4���{��������񚿒��i����Iy�����5q�i����&+	?-6u�"��i��V)���E�������X�iV�h��}�il��xJ�-B�#��s��Gc�����V�`�O����Ze/�4���>VDZ��+^��h��ʚ|�?��:0�����=���}B��D+�ɪ]C�Q�W��x�ŝ���!���8m���A� ��}�5,U����i��ʭ ��O�$ŷQi����U�Z��l�xF�ҳr���rcR����ZL�,�vF�簙
@�?LYK;䃬�h)�h0�9�r���	g>w�J�DVw� �;�)��폺���
o�Y߀0$F{)�9I�폺��"聊�� ?$g~ �t��Hea3r���u)x���
{�d��#0�9��u)0E��� ~H:��폲wI�C{�1XL�_ O\&�`$�J�"c�Q�YBk(�Ys�	�]�/�h��r���:b�R�6�A8�He ���B`z8LL�2"Ue+)U�8��VP�˙#d�p�GS�|)�Z���C
A�鋤R���2��t��)x�:b����LQ��`.2��;���Rb�� #|l����P\��^��Y��{�����Q�'+�������� ԰�o�I�H@鋤R�ĩc���a�:b��[��J�6>�۾�.%/�S&U����V0_,p?�%2��:b���q�X�|�����JeO�������X�X�Q�D<�Jf�m������1���dC��az����3XԱ�2�ޣ��y���!�\��;��u,q��w��"%3f�����a"
ǔ�V ��+	�x�0����O��ф�<~R9I�H��G�=X��E��{I�'���U �a'LU�I��`3X��E��yfœ�
?8�R�$鋈Rc���.���a����b��0�a��*A���1TJLt{�9�.���a+�yE�'�����&i#]Y��`$��M��I���c��1�	�1�(qYBk(�1�8@w��o݀0X��g��1�� hN?�@ $퐘�� ��7�̈�YGJ�Ue+)U�&��H�)�'��
}�m��^�d7zK���`S@(�԰��X���#�\e�-�wqv�6Do��4��w�H� ��B�O]�}�qo���a��_��4�i3H����V0_,p?�%2n��㻏������S&��������1���dC��L��Cw2����1���dC��L���L�V ��F��ta?m"̈́��a���.�i�q�@��X���M!ф��a��A̱wSM�R�����
h8�,&c����5|(�dA��_�ÃAHia3Z�}�b� �_�������&�	?�����]v�~�x(_�2Y�Y������Xt���P���o//�Mt�&iS;#RBl&���z�:���LH�� ��R� gI�c���A��H=�Ԧ@�y0�5֐��H5\G�@�x��aԒ�Ir��|�5g驁M����`@�8�Y�$&�q:A��eM4�c	Q0x�(��=ЎP==_R��W!��H8�n��C����$AQ}(0x�L�ܢ`����I�}/���%$>0�Z�_�/�JG�	#�}.���H�L� ��D<0x���LhnET_J:�f�}uf+	���!6���ͽ'�DǬ��e	��ʲ�=���A�Y�mfb����P	;d&'��� $��3"%VQҲ�YC��Ue	���6Jw	��u;�E�|�0�{"ڷ��.�k���MB@o�+�ſV��@�6Ґ.�kթa 7���߫I�A���?��yC�G�u�����a'�#�	{��en.��J�|���-̭��[���@��Y4�y�A���#�#���a'�#�݋^�Z��-K�o�+�ſr-D[���	 5� iV��S8V�4�)���!6G����C��ߙ�����ќ�����1M7�i1�$��R�Fr�<��B��39�Å��-Hu��&�xѨ+I�Huf+	��{�NDǬ����=�2n�����LŤ2�@I�!0	=&&o	�*������VR�(Mȇ�S�N#��>�-P��!�!N��4K��i3H67Do��ϯ4��~����1�vڸ5֬�W�GY�U��sY�YL�IIM���	a�lԐ��C�Hap�a��H]��s��' XoI��Hz�7��'+uf+	�����&�` ��O艏YG
�YI]e�{	����C�v~��E���)x���&b�@ $퐘�� ��7�̈�YGJ�Ue+)U�&��H�)�'��
}�m��{�R�M�����}����T��E�����(ũa p1+I�H|����q��l}��}�\_�L��m���݅����� ̈́�����	!��;em�v�Q�=�����a��4�o��� p1*�n`&iS;#RFa$s��}P�;�J۽��e� HI�)�)�I�5+�L!3��{�R�3���!儑η��{���S ~�4�NT���������f-!�N�	�@I��0	3xLȉU�t��VPⲕYBk.d����p!N���j��9)4�,��D�� 7��ۼJ}B@���kdC��+I�M[�>?t���b������ӏ��=�$s	?��ۨ���W�GY�U��s+0��;,X�7g��$w\��ң���Ml�x%V�-������	!�4v>�۾�.%B�=]�J�h�D[�2��э�E޹� ��V�4�)���9�$�p������%$0a$s�߻�䤄I�[��5�?���)]Y��`!�5�'	�c�R���T�v�ƈG����8�He ���B`z8LL�2"Ue+)U�8��VP�˙#d�p�GS�|)�Z���C
Iwy��4���w����n�u�>�l�!��6�*�.�_P�-��Gҍ���$.#ϻ��)�����n�Jff���O�����V�Y#�FʭD[�|�.��a0�f$&�`!�Ba0v����Bl&	oB����yVP��J�(Me=u�&���˘�OE�B�Mڿ������������3��'l���'��� $��3"%VQҲ���8��VP�˙#d�pGS�UO���rRh$�-��$t�����e�aw�_��Do�>� !OEZL�A�[ۄz����sH�a'�#��^���c�Do��LA�Uj"܏sH����a8�rlR)�g�{�S�1�����Z��$a$=6��Cx�)
lt i��)��17�E-���_1Ё���S�	on�3��b��LvC�a�&i?.��c������{���g�a0G��ӄ̈�j�YG
�c�P��k.o(M-��/B��G!�v���E8�� ��?�@ $퐘�� ��7�̈�YGJ�Ue+)U�&��H�)�'��
}�m�h��i\r�~���u�4��J������*)�(��jҢ�p�<�J�x��pwRKb��iQN��V�;�(�&i	�zJe����S.��a'�A��+���w��CK�6<�v���o�`V��Ÿ+�v���I�O\��	�R���˝: �;�#�՘�&/�J+�{�����L����L60	�M��A!?�Lz�<�(Me+(Me+(Me�\ǰ�r����;�A4��U��������z�p�&��YHYs�$8v���"Ј�He ���B`z8LL�2"Ue+)U�8��VP�˙#d�p�GS�|)�Z���C
K\K:^
$�n�H�Q�_P�]X��0�k�q�&i!����S04��~=����w\�� �,pah�p�9�-D[���˵� iV�K��p�o�FAo\T��_����@k��;;�u�p4[/�J�uI���OS�KƑ�3Y�a��+	�B����84Ȑ��i=pgd&=J�J�.t�$�4�7Vb����(���f�a0q�3�	��l`�0�	��:B����yVP��:VP��:VP��-���a�]�nA���A4ݸ�P����Dl`Z)�v�LOG	�@I��fDJ���e*�����Ys$l����w�>�T6��aI�!�)�'߀ѿ `���E����lg�a�Ȥ�j���_GI��5,$�8�X�i�,p7��ƭ&i�� E�5�X�q��M�IL��`�O�����b�:�*.�q}A�x�X��Z��+!�/������B@?�8;����l�����Q����7샫9V���O��z�M�+��J�T-��U��r6�e�*n��J໖�x�T/�ҳ�i��z���%�J�w\W�J��&iXI�iuc "���K�Cg����w,7����h��Ui3I뀓;!1�VRWYs�D'y�ź���E��Eox5Л	���|	��M��I�M��I�\&�` ����&=eU�&����&���&���P��-���a�]�nA���A-���4|]��!W`�������P	;d&'��� $��3"%VQҲ�YC��Ue	���6Jw	��u;�E�|�0�r^�TW��DG,
x`h��$wOs\)�v�oTzj%3sH2�����a7Q?�8��*)��j+�O�CK��E�'I��N�;�,ppk<\xz}�F6��UHn��t�hW��i4�I�M�a7��95�l�[y�p�-D[�M�=n��J��&i=pgd&=J�J�.t�$�4�wVb��	;C	��l`�0�����&����1�8Kh�4݀����O�V�}�Y�&vR@ $퐘�� ��7�̈�YGJ�Ue+)U�&��H�)�'��
}�m�r��((x�Q�k�`��(���f�����'��>��N����ZH|c���hH:��C�Y�-NHƁM�].dk͑�K5;< W�v�/T�e]Y�",e���-�ڴ��Ӑ���i#h���a���k�#�r�L��Ѩ`kJ��@����S>���M��zH�� E���f�#���S#��6#�S��"�z"5#��ԛ��)��*n@�z�0. �Sr��$8 �<����LvC��]"���S��%7 L�9Lyw]�
n@���C�-��ުLvC�\�E-#�S���jz���u�K�-�/l�U7 M�,Z#�8]z��p�;�A����Q}@jn� �����t�,ZG9M�c��z�Gx?�x*��'��g�#� �D�� �4��>6�S��bz:C(�� ����`f�B%VQҲ��ZUe	���6Jw�>�T6��aI��X`��HAm;"�h�v(-�Hia2�-&��/�4��®2��J�i�H��OU�4����,r�V����J�i�H�a:
���XjX�E-��J��`k�~��:G�������R?Yk�� ���&b��a;ncD��P�;R�'��@vݘ=��9�C��]�_�z�� �'m�w�E�L�1�Bnn�,;R�CS�����ƽ��S ���z�D�K-s��ف�	�wDspy%�߬��Α���|�?T��Z�I G+;nƐ�@ƈ=sp��v��=���D�ɐd���!w7]�TH�� Z����A� �"��sp��Aڔf��p �9�wDsp���o�Z��H��xھ ��#����G ����h����&�c�(��� ���r#�cD��7|OEڔ�v� C�vݍ!�"��z��=Cږ9۸�ʍ��&b�R=�(�nn4��ԣ4߻=  �E�6�	��4H����e��w� D�A9��4H����Jz�Q�p�1X)|�S!���Ɔ�jQ�Fvz F��V
���Bf)����cM��K-A�p1�Bf)�9�C�0v���vz Dp�!soi�S$sp���ݩe��;= !Bf+\��0��cD1���};R�Cvz G��!sob�S$sp���v��� �8 �a)��S!���ƃ7jQ�[�o�Z��H��xھ ��G�-p?�P !�"�/?u��4P1�Bnn�G�Ա�h]� %�f>�I��c@E$sp�	*v��KB�@~���1Yy��oz�E$&��	��Ա�h]� O�_��EA�E$sp��#�)�~�� r�(3�eUT�E$0sp�	c�/2o��`{� E`Gԝ�1�C�7p���.�J�����Pgo�h���� ɻR�%��`	��ڬ�E`B6�A?c$8sp�	h]�M(k�� 	��o ����л~��:G������~������f Gs��i'3ƈ=sp���K�����	��0	�v\�]3Ɖ	��Bhh�R�ӕvz F�(0R��S!���ƃ��K-�g�[�PgG�1Lh����!��K-�q�=s1Y��E$0sp�x;R���;�}��Ƒ���cD��P��K�������oކ5~�~�S ���z�D�K-]À�(:#��Gn߬��Α���| `�G�-p?�� F�"��Ҫ����cD��nڔҏK���f+8z��3Ɖ�!�t;R�O����EE���cD��n
nԪ�� a��	��i��4A뛀�ݩ�����9�?~6��cC�H�e����8��:O�o�"��)!h���� ��jQ�Z'c0^���"��X�4HA��OS�.�>.߬��Α���|��G�-p?������H&b�#���Q����9�?~6��i���\�`CUTA����؊Yiboz�f)����SCEڗA������z�#���cD��QH��e����Nf+!ʧm�h���$s�(�%N�4��3� �@ƈ=sp���(��� �����31Lh���'�(�ݜ��1XF� Nۘ� #��B��+�Wo�Z��H��xھ��G�-p?��?7O��PbȎ\"�����SNgj]4��  ~n Є��(:#��$���-ps�~�<m_ Y����\��-��V?Ҫ�s?h���'۵+�N�@ә��f� ��cD��n�jYi���fb��3lhL�1�Bnn�zjYh��� ����Ƒ�gm�h��7��,��;= Y���E
C�;ncD1����;R�M�ހ��y��Ez�o�l@��cD繸s�yڔ��� u����(E$sp����K����G��v4�w��4A뛀�9��\��v3  ��b��.!h��7�)]�t����Rf)�9�C���J3M��-ps�~�<m_ :���\�4 r���鋤R	��4C����ڔ�AހV"�.t�Y��f)�sp�����OP�� 1TJA3��1q
A3ƈcsp1��;R���;P "�DPa:�1Lh���!Mږ9-�������l�zh����%�v����o�Z��H��xھ `�G�-p?�=  h�Pe���oA�sp����K-�ٌ ��v������Yk��#���j��~������� �s�R	����.�"�����cGv��C����l`�����P1�<��HbnԦ��n� � Da�����AՈ�cD�n�v��M��f l`Z!p�4H��MڗA.���vݟ��"�����Կ��v� 60�����G*"��9�C��v����ܰc !����A7�Ɖ�!�v�9E"w� l`1��ϼ(�!���0M]�OQA�� ��.n"�!H�m�h�!��%�ڗA<v�e�t�߇�����R?Yk�� � ��"�#E��1�@G7�;�.���`c"~0B�E$sp�	o;R�'�;= ~.M���Pa�l@��cD��n=7jYiڀ�f+"<P1���i�Ա���8 �)3�#�"��z��=G�(�-]� r�(0R9�~�cD1���s�,d\��4�b�R`�4C���;v��G�gxOq�����yo�h�?Ϳ��4H1��C�ڕƋ�gxOq�&���[��y��E"����j�J�OS�L �����n4߬��Α���|��G�-p?�P �gm�{��P1�Bnn�x�K���p�EN����4H]��E�jQ�zq�pA���E$&��	�z�J3B����"��<�S$sp����R�E�c0���n�@ƈcsp1��v��O��=K�E����.=��cD��n�ԣ4ѻ� ��Eqs�4H`��=v�=KM�0 ���������-ps�~�<m_ ��#�����]�1XF%��1Lh���'(�K-6v�v��/�"��9�C�;R�'��4�_��V
FN�k ������cC�j^d5��@/�E^�s��4HM��C�jYi�;�_�C�En���cD�\� �1]�t�f��0	��m�B(��n�4Ժ��� \�"�0����f)�9�C��jS����`���.o3Ɖ� "t�R�#õ M# �����O� ���z��ږ9-��`2�۲�R�ۘ�!77M%NԺ	*v�~TEu��S$sp��ݩc��� b<�
 "���h���"�ڔ�"v3 �L�a����P1�@G7��ڗAgj ���L�cnd@ƈ=sp��ږ9���-ps�~�<m_ ��#����( o=ڄ�V6�b~��n�~�R�!����ـL�cw��v�ƈ=sp��v��� �Н�cw�D��4A뛀�jQ�[�����������P1�Bnn�uv��C�v3 ��"����4H����.��w������	�����\��W�p�R?Yk��&��s1XEͧm�h���'۵)�o�� .t���.���1�@G7�s�)�� ���n�N߬��Α���|��#����G [�k0����ә�cD��S�;R���;�]癊�.|�P1�@G7��ڗA=�� ��3�\���@Ɖ�!�[wjSJi;~��:G�����L?T��Z�H�w�{�'�sp��ev��LWj 3��co�E ���z�1ږ9n�^UUnf"�W�cD�� �y�ԣ4����\��W����~���C�&�:#���������(3/�`԰) ?-"mK��a�ҷL����&i ��H���`/ƕ�b<�Yn��&�J�s0���<�Yn��R.��}�W�oXjX4״�p+I��n��_�n�{r�i }ƈ��;)��԰Ғ �j�b�HR��r@����h)#i��L��*(�_P��#�L4fv���� '�G��,��B�B��ȩ�l�� i[���P��c@B9 �ߖ��J�HR�gF�!KM�fh��Z�����4�:a�}�	�>��L�� \^%<������O��l`�	 QKI��ٰ����4�:�J�H��c���X�L����95�x6(�l-�����踾r��r��'�����v�.����M�N�i3I�x��^з�������j�e,�yH+"� � �4}�+I�Nm���W{J�/�5�Yn۰���9�\����Q�s~�;"�2�"���H3 �4}�x�o- ����I�H��`�,��qo�4c��kc�}i#1h����_E}��kc����x���[��pkJ� ������ﰝ����jX6K��74�����/��s��a�mh)=�l0�3=�5�b�7:�6�h��F�� '�C�k� ����V�}��Ӥ���ƀ��>r|��yϻ_l��g��� k����/��6Q�wo��z��?4�6�>�� '�E�_F�ݿ�R�Iͦ����l�^�d԰�81�si�m�}3צ (��ZE��N�Aq|��u�Ɨ�m�w�H�1ƈ�bvRG_R���5,p7�� 5R���ZC�6��U���,T�[��I�\@ёu#��. ���^������ZEE��*-�+���R�׍IG�9 �c�#��������x7�>��Brr�O�i!67N�ɦ�o^�	�h�H<�8>��H��ct�V��X�$v����[l�ŏI��"�!p�Ծ�Ң�B����Ӵ���f���-l�?<'H
kVv�y�u�rԊ��4�V�����J��`k�� �z�H�w�G�"���X�iR=�e ͇\m\.4�*F0'�?
$3�0+IË�Rj+���ҭZ�5ֵ.�30��4�&��R�m|�5i\�A�,�8��k��JҤc~�� Q�F��g�/���C�;)��԰������X�!���$b�J�7�T^^���@԰������D*��C��5�q���b���f��Gn��Y)��큧�Wx��p�N�/�
�s`y]v���+:l1=��L��Dg�`_P^x�(��Ml�yH�Ң������K�A�H�Q���������'e&��5,)8[}��!���i���A�_��L{AHi�1�TX��a�J34�.�� ?q(�$m0�>�rrе炍�W���z�CL>�@0��`�Frw���Ӧߠ�|�%��e�i�l:G�?��೰�}�@O�����fc�}۰i��~V�}��Ӥri�{W��jDfz�n��a>��;�rrֹMK
T�=6�c�U�<8���/��@;T���u�_j�z�Bȁ��[-���^~i��"��x�i ����#}�a;)W�԰@m�i�_P�}V�K|�1��� ��R94ؾ�  ��,p`?i=�`F����k>�����7�x�V�K����#�L���!�C�ߖQ�_���9	�ڽ���"�M��:CJ��Ⱦ;@_�i}�اz���P��OS��,W�g'{,4��? �ԟ������������2��탍=��<�`X��ūH����l���ݚ4$t�Rm�+���������÷�Ëx�{e�}��!߁(���kaqx���$a9��y���G݂Y��_���� ���
?ge!��5,�ci�_Ph�ьC^�"�>��=?9V��ɦ���]��c��I��7ߧ��X��}  ''' 4Ѽ{Ģ��]6/��#i�����􀀜���A��ح"�M��:G&��'��C�>���,�`�->r�{-ZE.��t��0�����ol:ΣS���/ex@NN@#�)�t��6/��lѽ���:�Ҹ�r/�� ��Ƣڴ��P��OS��,W�g'{,4��? �ԟ������������2��탍=��<�`X��ūH����l���ݚ4$t�Rm�+���������÷�Ëx�{e�}��!߁(���kaqx���!�NECն:v�Ph�w�`�{���~+HE��
?ge'3��/Mό]��;{� iQ;����B��F�4���l�'xjX
>��m�����NU�r ��n!�d���In�U��\��b[ZC	ê����#����In�U��\��x=4�6�Ui ��� �vR���`f�ޥ��b{J�03V���#�G�A-'��i�}�z:v9v�N���4�y�{D�3q�藃N���4�}�t�P�ud�����}t:Ok�e����@Ӥ����5p����NHL}-�|] >���I�Ss4ٻN��(揼�����y1��Ӥ��<�!��+���t��	���OYҚ�\]��Ǵt��	���1�PP�ힻ�q5.S��>�i�{X"����2���2�r�CK������Â��}A�m��i�{3YA@>�;�.&J��p�Z��R�E�t��ZJ��H5������Zv�3I	�/�8Ԏ@	j���:��m+{KR��ft�(��86�����>
�@U�4����,�H|�|�y0�ZV��AP#�6�;���ґ_R��4��x.�6`x+I�CI���a�z�������ۦK""M�W��I��pi�����#�!I��A�ѻ
�iQKnj�Vo�� ��'�[�p�� k�(�C�^%��]jm��'楃KiR=��l�\�xQ����J�������6>� !w8,�sU��~���i!����Hd��r��`�'��h)�l]i�4�e�ɭ��������~�߁�,`:G&�Z`v��):l[�}��ȴ/�����6.��mf��f���\_9Gh����95�yZL�GoY)4����(\I���Y�<�楇�'��n�WNZV��E�nV������D���7��J����h�Rf�0�o/տ؃G�4�ҼwH��E\e��l�/��٣J�u��F ?��W.��_����h�i^��XH���Ҽj��ƈ�g�&aHD�,.��y~
�`(�����%%6�pY֒[WǢ�$@)��x�����F7�'I����E;�UZN`�#�0,�K�-*�[�w%�ȇ�f��@��o�ogxjX��P*a����������u,TS�U��'�������*C��`)�I
w઴�!1ƈ��3
C��jX
|RD��W�����F��5��K��5�K5V�4��iS����au' ��UZL�9 ��v�ŀ���.-�&�x�M`�,pO����#���qEu�v��������+I+��85�i � 1Ɗ癘RK�&��di[����}A�#U��'��'g�`��W�(�gPj��Q.����
�{p]*]BH�S����ҭ�B��v���n�X>�*)��l��l;aZ@� ����ﰙ�!�K�ѐ�d�$1U��Pv��:ݰ`V�A�V��}A�#|�Y�Y`V�h�v�>�|�?��DF13
H��jX7uƥ���$�X�#���+I�C⻉��Ԑ� ����.���7�K�+~�5��~ ��E�q��w
k�������ti�R��[�̸���]��R��Hu�T�ก� E#V�4�=�%#��l�2�c��H�05��6]q�p�Ҵ������(��`��$s/iI�4�����J�}j��ZԺH�8�w�Ґ��H}��եpil8������+J��	�+HQ1Ɖ~}�P��!��5,
6�ݰ4�Ӎi3IK�4d5QqE��om\y�}�_)�Ay� ��������o�N��5,#FF
���mZO��F7�`Y���vg ��h��դ� ~c}�{;�R�G�b�iU���B����RB�'R��#U��Ɖr�L��^5Ŏ���<��Q�5,`����t�����qJ�e�$v�,t����,�zȇ�!�+I�CM⻈�SG��431�`)�iV��kHi���2�4����*��%��������� �{U�b�v��}V�4�ۨ�}��l~. iR[���}�%$�]��G�ZBM��\�5���@��c=������4������;l>v:�K�Vc*����޲R0o�|�i[�Rj*'�IÂ��J�}��JM*&��R8�j�~0�x�i�O���"����i9�8���4���B��+1Ɖr\��&aI��������Ҕ�s��C�jX^<x4}԰��!�c*�u�X<�)
�흆V�&i/�F��?H�	�y��KN�J�>�h
>-+~�5��⻉{B/� ��Hy�j����S�Ҹ��f��z�H��X7��}��oiI�4��]$s�*���m)4���H�}�I�Om�Z>��6?4�-���>��w���#֭!&�V�o�c��� JY���_P�}�T^_��HR�;�v���+1�Z@���D@�3
B&@Ǹ��Ґ�����԰������E_ZT��MB�]��"��x�i3Hi�,:��~4��&�V�u���}��԰}����if1�I�G&�`���������5�yf��}��jX5���,�5i3Iz�H��XJ<jK�Vc/����x������]vH�Æ��v��1�~J�2��l8��i\��vjqv	I;�e��V�� ��D�(�A�3
B&�(�A����Ғ���R�U�<>��RF<,�xj�+1�P���U�a|dEڐm���H���0��'+|MK�9��<�I�H�y Q�W�J��d@Ҧ=a}D>
��]���dk}��E`V�V�o�/>�Bȁ�o�05��f��K�5pk�jX4oK���c����_)??ZV���
�ҷ����8R�V�4��JF�w���N@��_F����$>0��-�&�i ��cDa��>30�)_R��N@!���&i#u�F�_�*�͑J�l����CH��P�
����H|p�i4�O7��f�d@ҷ���i3Iͥ��5ֵ,7��JML1���J௔���+���}i[�A[�)�I�O��%#⻉{Cu' ����5F�M�+tӛ� 71Ɗ��aHD�R��zX�� _qc���πX�H7R�U��i3I��d�`�,7��JM:�Lw�X���I�Æ�&�ҭ�X}_�K�(Qf�+�i,8�����5���ҷ��R�_���Æ�d@*���Ҹ[�i ���E�(Qf�3
G%�5,��X��4���Mf����qk!A@�/���8�����~��� 5Y5�n���I�Iw�(���<�R�W.���p�ѩ@�`��[J�����J�o��S ?4# ��V��Ģ�����,.x�_�`k<�hȽ�dA�ZGMctڸ5ֵ,��;�/�q�Ĕ(�P�V�4��Ń^V���4c�8:�xt��i\e$.!�H8j�X��ʭ&iw��4��i���x4|�jM��6�_��<� ԰��)�5F>�i7 ��y:Y�{�?���{��Dx���r�����yK9aƥ���K�٨jX�i\���M��CR��{=�<+H �#p�J<j�f�J�����JC��԰h޴�
�(6�3T.��i�����o�I�}B@j�]�D+t�AZL�ȴ�u�|u,�԰�^݀���0+Hcm`f� � 1ƈ��3
M�jX5xW����GY�P�Wql�6�P���9;�a��8$�~YF�<i�I�O7��)�GY��h�iR"~�� � ����0�X�&��_��mZh�c׫I�E��čH� ?�Hrw��J^����>p^V�@ �
�m�덥n���8���K ?;�p�v���0%i ��Ɗ�,��P#}����!g'z��qc��!���԰���j+��$sH}�J�4�q���.D����!�K�DX��.o��s����\)?05�/ ��\����o��+��x|��1F�}cRr��u�����g`\J�~ ��Z>u,TKIu�q�<:�J�ҳ��Z��Iq���V���E����	�R<Md�n,p4�&��a�5,k��$����J��,fʬ�W�K"�t��+I�On�Pj�צ@j�:�5;>�������X�^��|a���7�i�4�U��{>�i � ���l�_3
G%�5,%m)u�@j��5�۶����Z����k��w:��9i�4�U�i)?�/���y��ʻ�xX�J��Z��#�3
O����X�iHa�5,��H+I�{u���8=2�/*z�)���m �1��I)�N��Z�F��R�wqL
�(5Q_ZTW��W� t���[JH+�J���I�CI�;��@�gR���U�%��{ 	m�� 1Ɗ晘R;�w8RsK����UdA�Ȥ��UB曝����m�4�:Nb����� ��<F6�������V������faI�!"�Ŏ������Wt��p�R�2���,���nhw���!���5�Y;	��*V�4��|���ni��.vڸjXp��9�iQ\e�	��1�|d�$>����'嚆v\}�|e,�x�7���RB�E�`��8�b��� ���!��mLB����|�U�FCU���ZCON��
6װj�[�{�l*<�-�HPJz����Ȥ��U@�Jo9��v��a��xp�W����)Ɗ��<��'5�.�#�Ŏ����`ѥN��\A���TX��� ��a݆���F��d@ё����Pj���ѐ�o�f�´��-��ҭW��. n��@D�����U�4��r�����,4��q����5!�Z�E�i[�Z�*)�����Ң[JEXp\^c�R�@��N�i U1�~����JCO�i3I�|I��R��4d5Y5	��-�!M��o�lg�J-��n��Q���F0ҭ;E���"� h�5��F ?��>-TW֕���X�A��� � �.J6�p=�0��|MK�\k}1_Z20UZL�~_��<�X�iH`i��["^��b�ą��e�� � �F��ȏ��3
B'�au�ҭTW{)��3�;,W��Hr�P��;�ci[�Vvĭ � �� �f���5,r��!��_�>դ)��!���
�A݅��ZH��uF"��N�J�r+�"��H���TKIZL�H(��l�y�]vk���m�%�� ��+�夃[�Z�4׈�� r ��#�!I�B���\M*-��RÌJE6���q��M�W���� 2�#�sY�&aHD�R��Kw�D<���ת�}��:OɌ,�xv��])������W��aԐ�U�q}@G^5&�	j���J�w
�h��;�i ��Bv�L��+�ܭ$`Cxt�vQ&�v*)ݩ`,a}��+�����8���� ���DF�f�J�,�Ҥ{G���H��l�$���B�M���ka�� (���0\^ ��k�A��/�P!޻�"�=��(�#�e�N~�����kaqHP>Ei3H��,���R�KTƴ�;�¾����i#�U-&��԰i^#���z��Î���
���oijX4�����]hRˋ���Hca�JC	j� ���"�3
H��԰�J��4��c*��H�0:�G!}B��t$-� <x�{`԰iQ_%�R<�����!��`-��\As�,~� iV�a}@Lf5$p�@�kJ�l��+�J��q�V�� z�i4���W���R��E��q�Fa�}A�x�ʅ�k�ҷ����WAI�᫃]hRˉZC��E�0�� ��E�\��a3
Nk�jX�W�\A 6���5
�s\|�o��*%��]E���oiY�"�����'`�r��J��+I�G%⻉{B/��=�ѨJ۾�x	`X��l�yI4�}�:�IZ@� ��
bD{0��|MK~4����0�
�������u��wIͿ-�K�֕�K�:��)e�DG�@�+t��Z@^ ��D��[ơ3
Om�5,�ҭqQF+�����Rc����S���"�Ml. �/�h��u�P���z��t��Se�^.ȇ�$A�~X}��$]�I����
�h5QN�5��#�uc���X��"�u�P԰iQtA}A�x�ʅ�3-�z5 � �1{��^5�$��ݼ�w���d@Ң�D>
����ö3�.u�\\��{@��Fҷ��,$m;"�l��x�XH�XjXw��ҷ�4~
�i^-5i ` ��!�o�7����SeB��� q�dC�!��T�&i1ȏDu��@� 1�D���P���Jf_OIq������Y�IY����-x]i�8�*5,[���$>5QN�;9��f���G^0� � �cEu�})�*H먵^Y�@_l�u�eXzT�o�Y���i��RXJ���&9莼`Ф� ��/�M�Hi{�6T/Mό_k�Ơ��u�"�o�E�-�"i����d�+"�J઴���"=׌:@M�#�
f!���u��.����v�$AgL��ہc���V걇5'��K	 ���Bgg`_Po��w`"��� ��U#b��%����o^Á�vv=��	� �T�#� ��U#h�(�g`<�ݴ@Ѿ�!Ŗ8'o��r ��A��6L��n ��3a��+��o���&���H���)LW��u��I� ~F�.��������RrM���aԊV�i�{���_�ȃ�aZCH�=���!m+;�lg����a D\K2����V�4��G�:�:�| F��ݰ��t�;��۷��@�� �Pf�Q&�8�噗+H���k����4���v���i3I�Dz#�) ���
��8|)gB�l�F�6�Y������Ԏ0�_�l�.�������Ң�E�p�{�8|)H�{h�|�Ų�
�㣵@E�$ �Gl�Yz�F@�F�'* ~>mWr�����4��c���#���~U����Pi����J��) ��iQF"���ZL�c�����@� ��Y���@
�p�H������;�u,7YH^���"���׍@R��@��ȁ�pUZL�<��Du� sR y���b<>�f:�M@��@���5#�� ��*�H�n��F9��t�JCK\T\�*&��8$�]�$�����
�}�H"��yP `�<
�s_|�����oTC���*&��&i��X�{B-�|���4��Ƽ
i��ZC-�iV��TM�ZL�c����M ��ch�&��q��U�A������au�Ң�_P����l��Ӫh�j�v}ECx��;��Nk�����;T�b-+rp�+I�G%��^ЊuVu������J�!��� 
�}�"Ҥ�*o���"���K3�["J��*Ņ��>���$A1�'�ʮ�׬��.�.+"J��+I�G�莼`�sH��ch�&��x��\�԰����⮬�20V�:�b�<�ݴAf� 
77N����ܫeZL�<����I� ~`G�����J�}
7I�Ipw�XM�A�H�Q���������Ŏ�E�iV�F�;	"��H�~�i3IYkdC��
74ci^`�00S;}#�����5��;���00;�;L�;�ݱ@֑�ь�q����j ��#��j�&���]�}�/hF��e���"��kVDEI���Pv��aq+I�G�莼`�.�������D���P��Rc�ʬ�4b�6�9i9��}��7ٲ iR�X�iD͢�t�RZT[y����q/��v=�H|� iR�Y�� �&��'��&��'�x5x]� �?)!v'G��-i��4��%!���00UUH�~��<5�xj%�"�	�⪪��� B|���UU#Q7Rf��Dz#�%�� � ��E|^n��u��v���n&Z�E��7���I��᭑R����q=7��6Tю@i��}Hi�܀.3n�u�>�m�81��E�Z���I1����&iDG�:�^� D���z��4p5ԑ���E��-�^�x4d4�j���Hrҷv#�T7�l�4���F�) ��iQF"���ZA��_��b,p5ྡx�_P�ūH� ~�Z�0xT/�ҤG6U�t���ٯ+��V�4�"#�x�,gH� �F����u�2�e
6>�9��h��,��|� ����X�������Iq��E��ȂH���	R�j;i
M��8��*|[n��i3H�"=׌�) k������B[ZCJ�H�z/ml�$�n���[jӪj�"�Hz"�z{�
6���Ѥi�n�P��0�����7�j�-��.��,Wi���ΙB������0��4�
��X��T�:�*.�	"7��S�#�OG�,ppR�x}j\ְ�*bRs�TQ�υ��RƤq�����M�N�԰<6�PV��m��WU��c�������K������ h��ZH�8�}T7^+��Ń_:���ȵ�w]�m�`1�r�8hȺ�ޣ��a��_�s �cD& �n�l:Mv^	�!��}�"-eZ���È�i3I���%�x���@�H� 2�>�W��
H먊f+���� �1^���w���ӤV� ���}A�E����Lp?���00L��"��ZE8��H� �vv1u,.hvk��i!�lf�;�-�U�� Ǎ�`#�!1_���j�AVuM+���M���kdC�� �9`S�@�=�/�#�'�ʬ�W��O���y���	f�@ �cEwF�\GRs=��*h�q��^5Ǜ;�;��8�X���+I�G�莼`=9�� ����pq)=�Qj��/ �C}��A_d^]!�N��p��5I��\L0���i3H�"=׌�:@� ����pq)#]�^^��E|���<��rwI��p��5I��\L0���ԑ��K�5p��sR�� ��tm+��B�	����԰iQ^Su�i �1���#�F��G��/KO��)G�F��N?zN�F2��J�o	��Rs1��4��W��1u,�@��i\?�aŝ��E�ޥ�J�򛭫I�c��iu�]�$]�ٮ�D<���O�_)#0�{�y��ܫ]��e�h�Ҥ�F�UHzÇ�a� �F��j�iV��aak��f��Dz#�c� 
�����yu��ZOm�^����]��@�#�F�&�ҸT|ۣ�N5$s��-�\B��D�a���8r�;���V�������8,���ZOk��-�g#�F�ga��o�(��qE���/��J���a���TE#V�a ��!�o�7����KeB��� q�dC�!��T�&iDG�:��B�Z 1��/�JI���Qo�;�5����a�8,�,�z0]������#Ȉ�G^0�R e ��Eu��B�F!�כ*�)�;"��+I�G�莼`=4� <��Es6�B/RF!���*�)�;"װ�+I�E	��5HۦԻ�k�j���!�ʪ���uw]�k8*�NӤ���� �})�;"�i%�����ͧV�p�5��9ZL�<��g�4i N���|G�Nm笰j���a��J�}
w
1:�_�P!اp�c�X�+���am��f��B�E�S�Q������+=�I��+�J�`_֥�Afrk�4��ġE�rk�p1RKG����&�18����ڭ&iDG�:�CB�� ��ݼ>�Q^�)Ǻ�sR�� _sO-�)W�\b+I�H�ZC�԰h޴��_�ž7LEڐl#�V�-�#D�8x�ӴZ����í�?��"�8Q���E�H�fȂJ@����O"���P\��)u٥H�*�ҷ�X���I�i�J��eZ���Ѵ���Ib��-*��(�_P� }/]���ݫI�G���c�� � ��#�G��V���.��G������p�RC�
�f��ol:ΣPn�J�|n����_�ZiQ7�NU��A���rp�+I�G�莼`��-����JG%�X�,B�IO��k�� G ��!N���S})��B�,y���*H¬H8������5��]j���3c��"m&�#H. ���|�BvD.����y����� � ���#|��Ng�#|l������R���`�^<�m)?��l��4�G�}������1U��0iR�ʅ4����R<
��?��+I�G�莼`�9�t ���ҋ]�E!@qH3{����Y]�������}ڒ�M��R�c�ZL�<��Du�t�@"�#
���(�X��b�r\`,p��[kb@l�����#�R�@��.(�c�Q��vv�~�;"� nl���g`[Ơ_PiV����o�w4h��ga-bg����(�a�d@Ҹ*�&iDG�:�8��v ��� ���}R^����e���ʚ�԰�8Ť�ۦ)LW�c��&i1ȏn��hR � �#h��q��#���!���z!���7��8Ť�n��1^���w��@�Rý�鴯���wH{ܦ�/ �����tڸ\�ZTNu$.(_�U��&9��x�
@���
����Ԥ7����Ǒb�	�F�4�����|X�!ŶT��@l\b�I���{7�ʛ����
>xR@�7�E �'����s���Sy�������p+��^�"��� #�_eM��qE<?�!6�Ja��������/�=K})��a��B��D)��ZL�<��Du�pΐ� �� Ѽ{ǥHi��X�;�Ѩ
1��T[xN_�A���D��,
u�*�C���_h�� \V���^=��V�V8��˛*k�R�H�_K�Ui3H�"=׌�Ԁ#����6T't��`C�,po�*o� 4l}dA%&�����4�����^��i3HzC�,po�1����*����$s}�T�q�.-�B"��񾈱|t�h��_�+�*���y����
@� ���t����u!�� ז8B�
�uMW���i��<��rv*��Y�+I�G�莼`���y �#
���Ԅc��iR?K���b����W�}2pg��@��p��  ��� Ѽ{�����<b�77�� �6ʬ�,^�-l3���ɩ`Ң���	 \V��=��gz��bJlggQ�k�?8�n� iR�	W�u����R�lX�kJ�w�&iDG�:�;��� ��|�?��RF����}B@h���Ȃ@!Ŗ8��J�%�X��鴫G�}���D�2��7a*V�4�"#�x�i�� Ǎ����ࠢ�CxYL�%֡�E�7�8��@���Ef���|����/�9�~/����<���IZL�<��Du���@~ �F>�^

 G���v�gq.�ŗ��*��VjX6F��ZNV疕R�濆+I�@� ���iE(�JIޠ+����-$s�@G־ʚi�H�n�MF�.)c���C� \["�;�o��x��ǁ�ZL�{w�	-�ؼ|8��?ZT��z��k���Ҽ?�E�1U��#Ȉ�G^0(� x ��|�?�1RF��G�F+"	 �|X�!ŶTѤ(۾�iI)�
R�ZV�4�"#�x���H� ��
�����Hz�b�7
S��YAAoX4������d��I�dC�CI�q[��[�M}�L��O�x��¿���tҼb�7��[�	��ZL�<��Du��ΐ� ��
�����H3�����\�����k��m)=��,p_��w]�z.k��8��w�H� ����,��p��r^!b��g���/J�1��!wv�#YH�/P�UCK�4d5[;��ȇ��A}���O�>���Y�~Y4����8����dR/��e���^n@�H���#Ȉ�G^0(~R �2�>k��m~Y�f���D8��"��]`���itĤ�߉�Q��x�u�x�1�8u������HR��j�w��� ѫI�M��'vmޠыR�x�k�g`э�H]O�m��5#���-J��԰iR�X� ͎��\����z�1��r��1�AP"� ��X
�i\%J�f�5⻈�P�K��F�iu�����R)p��W�R�����Hv ����4��y5p��sR��B��W���;�I	�S���gz�I�G�莼`P�� )�>�x�{o�k����R ��� �&�S��4�}��Bȁ�#\�0iQF���w��ʐ�*� iUv�!H
4W>D*C�z!𤀷�h�c/�k�/���n�.K��x��95���.Wi%���!�ۤ�v4O�iV�D+I��;/+I�B�x/�4�}�+g`��F�Ҿ�P�֩6D*@�Dl%J��a%������WHԚ �@��nTWY�v�A�h�(�LE�fht������@�_��j5��Q]a}u� i���)�����y���M � ��~l;������{h��z���I��t�jAm���tKR�@�D�%��z�3�,u$>jX]HH��/��f��Dz#�?i *��>��;����e�G��sR��vÛ�R��T����Ǜ;���h�Ġ����P�G�. iQX��붣��D<K薥�I�G&�a%����p4�
��ˋ�E�z�� �>1x������i]d}�G�)�VY�WX�^��I	�#�Y�J۽��Z@� ���Q���zm"�֓�u�(/X೰������ȁ�p��|�E��e�J����,w�'�$.;mGA�x����#Ȉ�G^0~K�i ��Q���c�e�$#�9�l��X(�{mv3�e��ޥ=`\A�ZE�1ZL�<��Du��� � �#(���Ӳ��ԟ�AJb�*)�/�4���P��O˘���B�� �1XX���f�"Rr������n>xb��� ���m&��#ƒ5�<��1u,?d�I��퀾�s_���(�]7N��W��1��DV�4�"#�x���H� ����l(�!����8gt�;�{OR��� ���yx���v"�[�ZCM⾊i��.+F9 ^^(/m݃Ȥ���"�t��#Ȉ�G^0~� ����MI��ź��:�AE�u�H�cw�;m�'/�,p\mť�`V��.�7�4i"���`԰}�/�3.(�3����o�ZU�����ܭ&i=�QJ�8��[�iQqp�2kaqRs5p�ȁ�Z>��Y�ph5�x5���I��(�u�K�$�(
7_�@��PP�1쐢�n�i3I��X븗�"�V�������d���i���
���"N�+�>1U��#Ȉ�G^0~GR � ���!I��q��^Y�$�&7x��r����Z^i9��&��#�R>�l��4�G�~��f��Dz#�?) � S�,|B��}ⴊ.�#�R>�l��4�G��j���ȩ?TQ�π��!��x+sȟ����+s��`'�0n�W����$&�膱Z@)��
���05ԃ;����-�h�ly���[�	�!��M��/�}�}_ ��ѿ ���wv[��7!�i�-�װk��m��@�ZL�K!rҭ:���FF
����
�h�V���m�pUu�5/]v^�y5�`k�����y�-�'秿��`�E�^xdC���MB@�xjf��)�\���t�p��
��̸��'�"+HF8��X�l/Do�Φ�O�= ���Ke�i��sZ�T�'+|F�{s����=��F7�m�w����Ҁҷ\W�m�Ҹ*�'�������K������ h��ZCK	�}T7^+��Ń_:���ȵ�w]�m�`1�XKFE��&����� )FѴ�*� ���uqZ�^�԰Ҹ�i��qc�o�'�|h�ҭ�\ʅ�$�8)85,06��Q�����xu�4d�d@"+H��#Dmn�stHS��ZH�c}�t��*���5p���t�F�]�a�X�5�!�`V����}A�E�. ��T\[�6EI௃W���Z�A}��
$}(�8|������9볽�Rs ��i�gxjX�_�*(����{E�ÂJNf�/�m�b�7
��Ku��EŲ ��V�� ~c}�{;�R��KJ��xIn�!�q�I�	���Ph�]q�p�ִ�����4�է�2��`�5���=��p���(�["����i[���n�u�l۰�N�3W�֥��ZU��_ZW��O�5'��#�6�;�R�U�+��ZG������K�-*��F��\^F�[��x~Rx�d�,�4�\m\.u�*'� �#EjQ$G��Ez5ԟ�×��A�A�o���C��St��RZy��iQw�;��V�SX�_��H��p�5,%5	� )�yF������).���.���V� )�(����;��P��� ������$C�\QzERŵ�a�s�k�c�^�^�����{�P�u	�Ƥ� ?1��:N�԰l�+�/�(;n�n�!�`2)L$C[V������w�������9x25�i4 ��o�ogxjX��P*'��m%�ȇ���$_�;5�%�W�k_?ei �S�+��/�����A�ZG���" �������J�Y��/�j]"�~�ʛ�gadA 4����R{ZTQ��ժ�㳰���(�������#��`�"�m�4��]@O�ZL�8���Q W-�Z|M<�>8�q��`k�w���֕��#�	�R~jX4׷�
�s��U�t�<�H� 1ƋSc;:�C�����\�}�اxYH�n|7�V��}C���n|��l��|Y S�X�i�Q�ȩ�*�����w:�i�)�=j� � �F���}�a�Z�'������jC������_v"��i^���(#��].ub�\�Ԁ�GR��E>\8���� ��0,���Iu7ߧ��Ph�s�ѤۦSQ�4o�p�%$q��B�O�P#ҷ�����Hd�-vG֚7\f{���ȇ��6�;դ� ��:I���z8�T�]�x(^^�qU������ �{I�95�߶ڵp����t�yZ@{ ���.�B�^��_����v.�B�7������ �PiV��mZU������� �Ɗ��>8bRh^&�*)�n��o�Oړ�Q��P��@����O6E޻H�� � ��"��͵�jB1ŉ��K����J@V
vq��Hy�P���n^X�c��04o٨Y�p7/�ei3I�C��J������������xa&�qRl��$Yd@ҽJ�����<��4��lS�Z@9��y��"�CM��\�@_I�w�WXHi�G����,�/��v�F�m+u�&��v�'௭*A@���s�FG�]M��P0���ږeH8V����T�����Q�R�����>�O��P���28�V����z���05ԑ����x���/�,�|	�x.� O�E�Z�>ECxp�:K^���ȇ�ё|c]I��Rۧh��$�8��R~ �_@m�\[�� iR�%K�� #!#�ZA���T���Y/�jX]I�H3a���PQ�'M�a}����F�ϻK�����Î��m�m�_|V�� ~|Nu�}��7��E޻H���)0�� �$}(�`_a����ZC���4�}"v�P�0�-�r���(Qg{���9a�FF�vx*��n3�*�!����԰�-zΣPiV��Wȭ!� �D��h�췁�{ ������m�=�P9��ÌG�=��Gl�,�5,�Ml. /�H��f���c>ܮ�Z@� 2ƈ�Z��F����v��
J��u��28>K���qM""��|��(���U��P�.�dC�i���ҷu��,pM����i � ���;Mu��'��-x/�4���O"�DE�a��I�QgM������O-�>�Az�u��D<5ƒ5Haⴀ� ���1��򐁰����Á���m��vդ��^�-l�fû����6>�w�����aԐ!��frr+H7��E�F��io�7ِ.|��g`+�ѣ� �*B��>m���f ~{���W}ƐU'�����y0������C���i�U��^юJNf*���`+�q���{c�9#RC�	W�7��G���%i � <��o���c7��G���
T��/m�u�a݅�P���f������c���&i^Q�Uu�W��ȁ�_�I�,pY_sO<.�i _F�o��1<0���B��a����S���fȣR ��"���	F�+���i4 ��"���	"WVD�`W�i< ?��7�$���'a%!M��h�p�1���&i4&��o��6>w�ĸ�a���w�Y�Y�'�v�e�����x� a������dU''a 4�>���iII�c�.���X�r�6��,-x,�������j�f[�B�]q4d�,?zl>켰g'{R~Yz�"�E��7����f�~��j��{�����}�̾���e��-v�Ei ����/ϲ�����fe��l}�r.v��D�t٬��\]�}B�,W>=��{l��򴙤��i���/<�!�
?�n���Ml./�-�b.ԑ½4Z1�w�v���n�B�H8kHi����=��HQ���߭�.�!���>���԰�ڪ;��;����EŶ��_ZEm��}2�ɮ�������r4~���9ZL���C�:e
,�5�!�
0,p�����.�m��V��������#��7ِ��gadRJJ.Pu�k�
���$c2�h�d@ѧf�ga���i���])��R9���WK��<��4K�5�=�)#vXj� ]Jd����ܨ=�ۅ��4��N�Π����eŨ��3Ա�P��*Z|syI�� U|a�]�C\Q����J�[",7�(ŸW����ONM����y�
I_�� ���҉�F ��9�"hъ?��s�o��aw�@kթa%$0o�7��f����a����-K� �{��R,�HԐk���a��>դ�������;(�����i?�~0��ҷ��� ��(���g�����6>�p1ŭ�kaq+I�O��a{E�a 7�.7�G�Om�(�L�� 7Qt}�:ȇ� �Yq������q�ڴ�� X�/��������
G��^�V$ʛ�ga��I�ȃ��+��Z|sx~�n�'������?r=���v蹮�*Ha��X�uդ� S�/�������|i�AzEX�*n���E!��u��`W��X�#�``/+H� R��� w�7��,p�00�P��eVv�5�}Ŏ	�4�V�K{��5i � Ѝ�/��n���M'1�EP>�/�A�o�u��E�IH<�J��c �!7?�|[�����|i4�6Ug`-��@�� S ���y�=��Oސ�����a{|G��i 7���_�mӴZ��G�c��=K��"WM�j�,\=�¸5u'`�r�����X���Z����E��7�gPj�+�����N����9��_�k��m\/i�X4~��c���IrD���C�%���çn��y�=e�/���H9Z@� ���(�G�`�����[F��m���p�_��V�4���oj�V��� _��V�Rƈ��ޠ����QqJ�wR{t���!��� �UUH�̸��s����C}��Ha�	�I�F�C ��*�}���5	 S�Q����V�4�M(�Nz��F�癗z�x3׿ �������JOv�
��F� 
w
188��� � �0�7}Ŏ5!��}�y�Ԝ׊��]K	�����*+�� ���ʡx�u�R���`ҽ2Y
|�I�/�s_}ŎK	��_B_P�V�_ �#E{V�Dj%�"��vk{Vʮh�c���a*V�` �#
�w�o�%�$�ö;�ڶUsE���kH6�T� � S���Y^�KH�6��jG݅�����\�#ǰ��s\'��Si[���ok��� � ��¼�M{F5���uIx�쩌�N��E�i������}Ŏ	)�|Zy,p6>�nV�4��1���]�I���d�T]�o��h��I$=����� �#Dm�kaqw�e!�]�b�X
|\>��ɩ~�qp�M¼����4��884U�� ��DR:m������2]E�� t����,�Nr������q��}���5	 H�P"���CK�z����Ң�� �%�a9ѩ3H=��M)1�@J@��"<蹮. !�$x�F�R�O���Q��aqv�1��X/l��<���������z*�⾊o�)?/m�T]�ʬ�T����c���#[��+I�G&�`�����$9ꪩߞ�SF6����/�IIKi�4����. i[���wY'�FF
�_��Gſ���z�}C���eXZ���)ƈ���x���c��>���P��/�4��jA���6�
1�jl�W�J�}am��f&��$p�=�k��2�����J��}B@�N���|h� jl���LE�f5�Xa-�jX/l Գ95�V�������@B�#�l��b�U��EI0��vp� ��ƈ��ޠ��7t����#eE�	 �Q��N���"�4�	R�C��dr��xu�4$���A�u�s�,l=A젠&��9o�u�X�L���W�z5&i,&nF\��>V�|�g�`�R)XL��h�:E+	�(��)0��%� ̈́�j�+���$~��H��攀@�#
�zC o�jPY��C
G%�t� -��6����UU!����Ë@�&i#-��w(ט�&ҺCUVo����j��M��u�泂���:A������i�����Ɲ�o�J��ÃH`����{~(��� a �#EjPY��C o�F�C
E�e,�",/o��H`D����UUhR��+Hx��#��ZC
M����7��R����ZNlB�v���|�����}��\�E�z�C
L|=i3I�n7�K�F�Ʃ6��*��x�P����T��m4;��5�T'i����$��]��H`����4�xx��КT��vCUT����G�|8�V�h ��H�CT�ޕUVoU"��@G�C��U��}���$	�*��ުA��i d �cDG�l�Rj&ʪ��JA��@G�l�Y�7�k�}B@Q6UUf�R��+H\ ��Q6�Sq)1���i��h}�M�UY���l%J� <��!�o��mH3����`k�x����C��U�����Ԇ2��ZL�H�xԻ�k�j�iUeUVn%$f�]�ڤm�i��v��ડ;N���7�$A�0���RvD<4,
�M�URF�X�ƾG+Hp )Ɗ���Dj'>���O�ߞ)�u�[@+씐m��?�+H_���!��HN}$k�ߞC�S_dC��/�!�����u�[@X��q+I�G!�o�y�Rm*'=UU#Q9���uw�j��M��u�泂���:H�sxDC ��o� q�dC�#]!�
hX���UUH����X�ƾG+Hp)����o�'>��u���b��/�!�����u�[@X��q+I�G��o�r�y�Rx���������:���Hۦ�Cv�P��ઠE��7�$A�0���RRxӲ!����4&��������]$x�È�i  2ƈaa�e�}��<[����)��@��X�i�'a q�!@a+�K	��>8U�a<ƈLU�l|+�s]dA��ICW`_P�0�k�_k�}��5�'t���U->9�����(;n�����W�#���@�Ѭ
�|c/������5�e�ԙ�������{���I�Om���7�{[��JI�a��/�HZ5�\/�`��Bvz>���jL�@R{(��ɹ������(�Hc ���#ݾ��ޑɼ,���E�����dA t�kb��wt��� � �#D��t�;k��k�í�^���>-<�W|a�X�>�G �m+|a�Y}A�H�0�.�ʋIZV��%J� � 2F��/-�. xA�I�{����W���w6���� ^<ln7R���� 	*� ��D���1)#������1�=�������K����7LH�V�4��.�Ң�\d�$����=� ���!�kvÆ���3W�!> �? ��C�	U$st��԰n�c�]qb� {�#�Z@� S�/�Ν���z4����اw����+ц6k���'��2_�C��m*.��%J�f��r_ON�k�_�[*�iII�c�to�u�:l�]���� �#D`�Ӱ�����Ne�F�;E�`_P�~��+�s]'`'�I��`%��&i?�(�vt�l]���H:�J6X�i�&�Ip��.�a�M���u ���p/�^�KI�u1WOx�����;0�]v^T�T���h������K~� ] �F��\C�b/�q�'�� ��х��J�c��x�E�0V�� <ƈ�q��
�\�Y]�a��8�� �|�]v���5�e�Єr����[���iUQ���Gw��>o�i #)F���X�����"�'5��
uM�*�������̝�i.1�Ud@(�7�UU!�l��vDR(E�z�zUUR�ʅ4&��˕ 0۽v^�P�Ҫ���7��h�^��Q�E�5w�����
�8.1��HM �F������E���<�x�Z5�\/�5˾���g���5���A@�?�ED�C�C;B%BB.G�F�F�J�JkJ<J�IHPK?K)KKUUZU VBf�fu��ńQ�|����+������n�r���%�ڌgg!gh�	h�h��                                                                                        [mouse]
MouseType=Serial1
>>  R6000
- stack overflow
  R6003
- integer divide by 0
 	 R6009
- not enough space for environment
 � 
 � run-time error   R6002
- floating point not loaded
  R6001
- null pointer assignment
 ���                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 ; SCANDISK.INI
;
; This file contains settings you can use to customize the ScanDisk program.


; -------------------------------------------------------------------
; The [ENVIRONMENT] section contains the following settings, which
; determine general aspects of ScanDisk's behavior:
;
; Display      Configures ScanDisk to run with a particular type of
;              display. The default display type is Auto (ScanDisk
;              adjusts to the current display).
;
; Mouse        Enables or disables mouse support. The default value is On.
;
; ScanTimeOut  Determines whether ScanDisk should detect disk timeouts
;              while performing a surface scan. The default value is Off.
;
; NumPasses    Determines how many times ScanDisk should check each
;              cluster during a surface scan. The default value is 1.
;
; LabelCheck   Determines whether ScanDisk should check volume labels
;              for invalid characters. The default is Off.
;
; LfnCheck     Enables support for long filenames. The default value is On.
;              If LfnCheck is On, ScanDisk leaves any long filenames
;              unchanged. If LfnCheck is Off, ScanDisk validates
;              all filenames, including long filenames, to ensure that 
;              they conform to the "8.3" file-naming convention used by 
;              MS-DOS versions 6.22 and earlier. 
;

[ENVIRONMENT]
   Display     = Auto   ; Auto, Mono, Color, Off
   Mouse       = On     ; On, Off
   ScanTimeOut = Off    ; On, Off
   NumPasses   = 1      ; 1 through 65,535 (anything over 10 is slow)
   LabelCheck  = Off    ; On, Off
   LfnCheck    = On     ; On, Off

; -------------------------------------------------------------------
; The [CUSTOM] section determines ScanDisk's behavior when ScanDisk is
; started with the /CUSTOM switch. You can adjust these settings to
; create a customized "version" of ScanDisk. This can be especially
; useful for running ScanDisk from a batch file. The [CUSTOM] settings are:
;
; DriveSummary  Determines whether ScanDisk displays full-screen
;               summary information after checking each drive.
;               The default is Auto (ScanDisk displays the summary
;               only if it encounters errors on that drive).
;
; AllSummary    Determines whether ScanDisk displays full-screen
;               summary information after checking all drives.
;               The default is Auto (ScanDisk displays the summary
;               only if it encounters errors on any drive).
;
; Surface       Determines whether ScanDisk will perform a surface scan:
;                  Never    (Default) Does not perform a surface scan.
;                  Always   Performs a surface scan without prompting first.
;                  Prompt   Prompts before performing a surface scan.
;               The /SURFACE command-line switch overrides this setting.
;
; CheckHost     Determines whether ScanDisk will first check a host drive
;               before checking any compressed drives located on that drive.
;                  Never    (Default) Does not check the host drive.
;                  Always   Checks the host drive without prompting first.
;                  Prompt   Prompts before checking the host drive.
;
; SaveLog       Determines what ScanDisk does with the repair log file:
;                  Off        (Default) Does not save the repair log.
;                  Append     Appends the log to the previous log, if any.
;                  Overwrite  Replaces the previous log with the new log.
;
; Undo          Determines whether ScanDisk creates an Undo floppy disk.
;               The default is Never (ScanDisk does not create an Undo disk).
;               The Prompt value causes ScanDisk to prompt you for a disk.

[CUSTOM]
   DriveSummary  = Auto         ; Auto, On, Off
   AllSummary    = Auto         ; Auto, On, Off
   Surface       = Never        ; Never, Always, Prompt
   CheckHost     = Never        ; Never, Always, Prompt
   SaveLog       = Off          ; Off, Append, Overwrite
   Undo          = Prompt       ; Prompt, Never

; The following settings determine the corrective action ScanDisk will
; take if it was started with the /CUSTOM switch and finds a disk error.

; The next five settings accept any of the following values:
;    Prompt     Causes ScanDisk to prompt you before fixing this problem.
;    Fix        Causes ScanDisk to fix the problem without prompting you.
;    Quit       Causes ScanDisk to terminate if it encounters this problem.

   DS_Header     = Prompt       ; Damaged compressed volume file header
   FAT_Media     = Prompt       ; Missing or invalid FAT media byte
   Okay_Entries  = Prompt       ; Damaged, but repairable, directories/files
   Bad_Chain     = Prompt       ; Files or directories which should be truncated
   Crosslinks    = Prompt       ; FAT-level crosslinks


; The next seven settings accept any of the following values:
;    Prompt     Causes ScanDisk to prompt you before fixing this problem.
;    Fix        Causes ScanDisk to fix the problem without prompting you.
;    Quit       Causes ScanDisk to terminate if it encounters this problem.
;    Skip       Causes ScanDisk to skip fixing this problem, but continue
;               checking the disk.

   Boot_Sector   = Prompt       ; Damaged boot sector on compressed drive
   Invalid_MDFAT = Prompt       ; Invalid MDFAT entries
   DS_Crosslinks = Prompt       ; Internal (MDFAT-level) crosslinks
   DS_LostClust  = Prompt       ; Internal lost clusters
   DS_Signatures = Prompt       ; Missing compressed volume file signatures
   Mismatch_FAT  = Prompt       ; Mismatched FATs on non-compressed drives
   Bad_Clusters  = Prompt       ; Physical damage or decompression errors


; The next setting accepts any of the following values:
;
;    Prompt     Causes ScanDisk to prompt you before fixing this problem.
;    Delete     Causes ScanDisk to delete the damaged directory entries
;               without prompting you first.
;    Quit       Causes ScanDisk to terminate if it encounters this problem.

   Bad_Entries   = Prompt       ; Damaged and irrepairable directories or files


; The next setting accepts any of the following values:
;
;    Prompt     Causes ScanDisk to prompt you before fixing this problem.
;    Save       Causes ScanDisk to save the lost clusters as files in the
;               root directory without prompting you first.
;    Delete     Causes ScanDisk to delete the contents of the lost clusters
;               without prompting you first.
;    Quit       Causes ScanDisk to terminate if it encounters this problem.
;    Skip       Causes ScanDisk to skip fixing this problem, but continue
;               checking the disk.

   LostClust     = Prompt       ; Lost clusters
e o � � =d��0&'*u)E)((�'�''�&�&�+�+�*{*�+�+�+�+	,,S0�; 	0&x0i11�1#33�3w4�8 |<`$0&                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           ���� � ! MS$MOUSE    .� .� ˜S.� �w � uPQRWVU�6G]^_ZYX��G ��G�[��      @ ` � � � �  @�� @�� @�            ����  ����  ����  ����                                                bc � @  2      22    �� �   P  @                                           � em                   ��������������������������������                                                   �    ��n � �, 	�)��G 4� �
   �+�  0 ������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                  �?������  ?  ���0���   @ ` p x | ~ � | l F      � ��� w                            �         � �   ����     �
        �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              !   8"8%((2_�����x�)�"37=CV���`f\<��$9JQ�� 1cx���`��^��	
 !"#$&0@t~@ABCDE`ab`anopqrxyz{        		%')+	!%).	#'+05< $(,0 $(,048<@ $(,048<@DHLPTX\`                                                                                                                                                                                                                                                                                                                                                                                                    *** This is Copyright 1983-1990 Microsoft ***��8.�� .�� <.t
�u��.�� .�� �.�>x
 t�.�� .�� .�.v
.�� .�� U��W�v��v
��v��v�<+t1<.t-<	t9<t-<t1<t%<t)<t%<t<u!��T�|�t��������t����ߎ�P��~��~
��~��~�X<,t<-t<t<t<)u�~
���~��~�5��v�_].�� .�� � .�>� tx�Ȏء@�>x t���лs�?r
�?t�?u����=�v���>� �СB���>� � v���>� ���&� ����t������� �� π�t���u<0u1.�� .�� .�.r
.�� .�� .�>: t�r
�u�.8&tu�P�� .�� �X�.�� �.�r
.�� PSQRVWU�.�>; t	�ˎ��+0�13��ؠI$�ˎۻs��8&:t
P�F�<Xr
�~t:t��)�#�����E]_^ZY[X.�� .�� �<2s/PSQRWVU���<.u��2�S����،Ȏ؋��
[��]^_ZY[X�<Mu�ώǿ��<mu�ώǿ���F �7���9 w�s�>t u<�>5u�� �-�>; t�\/�'��� ��� $�>5u��P�Xt�0�s�d�2��;�>9 t��,�	��  ��  �� H�� �� H�� 3��q�r�� �� �l
� �ώǿ� �� �D�F�wH�� 8~
u��������0 ��!�>9 t�*�,�f����x����� �� �����s��3��ؠV�ʎ�<@t
<t��ð#ð&�;�|�ʀ>x t�������� �� �>9 t��(�;�|�ʉ� �� �>9 t�(��� �� �����؋������ �� �>; t�>u�>x t$$�� �>; t��>�.�>; u	�>x t$��@�À>; t�>t�>; t	��>�.�B�>9 t�?,3��<�>�8� u�Ȏ��q�N�q�����،Ȏ��� �n �	�	�,�	���)�	�4�G�	��
��~	��+��v	&89t��9�[�g	��Ȏ�3��289t�)�+3�넻� ��?�u����� 2�F8&x�@t$��F�B��F
þ� �t�� 3�8x���F�Dt$��F�D�F
�� ��Fþ� �tվ� �Ѐ>9 t�h+���� ���Ǌ�����>��.�����F��Ø�>; t�>u���t�����D��Î��=�Ȏ����F���2��� 8� t�>� �u�Ȏ��q���q�� �2�89ua�� �;8;t�u��2��+�+��t8Rt���� w�7�9���u
�t@w�t��� �"�"Ԋ�ʴ�� ��� �3���� �F3��� ��F
������� ��uA�uB�� �� À>x t�>; u������������ �� �6� �>� � �� 8.� u���B�@�8t8.;u�8.;u���� J��� I�28.;t8.>u�+F+D8.xt����BB������JӋ�_I�s�>9 t��)�q���q���@�B+S+U��t��� �~��� �F
�� �F �� 2�F��� �� ���� ��>�  �u&�> Gu
�l
�!$��!��Fk������ �n ��	�,����)��4�G���
��|��+��t��9�[�l�Ë��mu��F
��F��F�3��F�F
�FH�Fød ;�r��;�r��;�r�Ћ�
��¢� ���� �â� ���� �Ƣ� ���� 3��� �� À��� �>�u�3��� �F�� �F�� �F
Ëãi�&ge�cái�F���5�~
�� �!�� ����;�u=��hu7�r
�t
�>� u�>5u��4��4�ظ%.�� �!.�� �Ȏ��r
  �j
�5�� �!�� ����;�u*;�u$�j
�%�� �z
�!�Ȏ��� �z
  �>r
 t�F���x
�F �v
�FÃ>r
 uj�5�� �!�� ����;�u��htO�>5u0�>� u��4��4��6��ڋӸ%R.�� �!�Ȏ��� [�r
�t
�%�h�� �!�� �>z
 u8�j
�5�� �!�� ����;�u;�t�z
�|
���%�j
�� �!�� �>�u�ˎۻC�� �� ·��� �/ �3�F�t�~
 �#��3��F �7���9 w3���;H�F�>9 t�%����w�� á� �Fá����F�����Fà� �2�8&;t�>u �F�q�F�� ���F�� ���F
�2�~
�F�� �F�� �F
�3���� �F3��� ��F
�7�F�9�F��'���0 ��
:tC��É�F �t< u2��s�[��t�s ��u�u�
�u2���u�N3��F
�F áD�F�F�F2䠟�F
�� �F��F���ǀ�s؊�2��࿈
��%�R�F  ÈQ�F  Ë���r���u�����D�L�D ���F��Ã��u�,�F Ã�wBK�����،Ȏ��n�� �Ȏ؈$�'r�%�� �)��'%��n�#��N��F���3��F�$@�F�N �Fn�3ɠ$���t3K�����w*���$�'r�%�� ��'%��n�#�Ý3�2�@�FH�N��������r�N �FÀ>) u)���،Ȏ��  �r���
�t	��.� �Ȏ��F  ��F��À>h
t�h
�F��h
 �>�u�6�FF��s�F  À>�u��>�u�� P�� P�m
��2��� � � � JJ�j
�5�� �!�� ����;�u;�t�z
�|
�j
���%�� �!�� �m
������ � JJ2��� � J�`�� � ����� � B��� � ����3Ɏيl�� � :lt��E�� � :lu������ � ���R�� �:lu��Ɏ�YZ�� � ���� � ��� � ��� � �� t�>� ��� �� u�
��F  X�� X�� Ëm
����2�8�t�@
� 

B�>� u�>�tJ�G��������u�2PS3�
�t<dr�d�@@���2�X ��؋[Xt�2 ���s���Q3����"�t"� �� ���D"�u��:���uY��t��Y���Yó�B�M.�m
����3Ɏ��+ �u
:lu��������:�t��u����Êl.� Êl.� ÌȎ����*�n�� �"�$���'r�%�� �&$'%2���n�#�>)�À>�uS� ��� ��� [Ë�
���� � �k
��
��À>�t��
���� � "k
�À��u<v<4w<3s<1s<$w<!r���Ð��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������s�{����u�� � � �x� � 3�8qu�8Qt8� u�P�P:QrɈ&P�� �>9 t��tM������<Ù�>� �<� ���� �����t�>; t�>t�>; t�����@+S���F������>���>� �>� ��� ����t�>; t�>; t�����B+U�Ȁ>�t�>�t	� R��
�Z�� 
�t52�8&ru-�rP�� $�t#��uXP#Dt�D�u�DV���� ^�L��:XP"� t�>l
 t�!�u�� �� X�t��� 
qu��q���q�r]^_ZY[X.�� .�� ϋÌʎ��G >%2��R���.� ����� ��׿ ���� �؋�Z���.� ����� ��׿ ���� ����PQ���y���y��;�s���>'2�#�O�s���I��YX��3���&�$t��s�����Ȣ� �2��� �@8>xt����B�6� �>� �� �>�^ �.�� �Ȏ���Ìˎ�&�>; u� ������H 3�&�4�`�; &8;t����+M� +͸���͸��� �� �&��AA��;�r�&�_�.�.���.��.�>� u.�&�
�խ��Ju�.�>; t�ë��ê���V.��H.�&��؋Ȭ"@�u��.��^Ëխ��3ëJu�2������

��ϋ5���B���J��B�����Ȏ����>9 t�+�B�@��}�{�>ty�>; t� �>8.;te�>; u��� �}�{��� J��� I��	r@;� s:;� s4�	�>6 t�5���u���t�&�����2#739� �}À>; u+D�>x t���H+F�J�>; t�-r^�>> t���E�>����7��BB������JӋ�_I�Y	r)�X��N�>st��;�O� �{�S�}�U�2��28;t�}8t��>t\8;uޡU�S���2�8wt86t��5���u���t������G86t��5���u���t�����Ȏ����d3�8	t�8;u�
��=s��8;uG�3� ��ں������ � B���J�ĸ����� � B���J�Ĳĸ���� � B���J�Ċ����2�������������}	��� �� ���߹ � ��߃��� ��� À>2 t�W��o � �W��o��H�6J�C�����`�.���>; t�� �&�
�؎��խ#3�CCJu��"2�CGG��Îy�խ&#3�CCJu��&"2�CGG��Îy����&.����>� u5��BU��&�%����&�%�G�CCMu�]��&�%��CGG�۰��J��&.�ð�BU��&��&���&�����&��&���&��G�CCMu�]��&��&���&���CGG�뫎y��S�?��� [CFJu��>; tCF�����&���r2���s4���u�Ë.���H"�"4�4*�t*|G����� �Ǿ`<s�؋����G������Ȉ��u��V�َ��ȋ���2�2���
ÊܪJu�^��؊���� �Ǿ`���N<s�����O����������u���V�َ��ȋ���2�2���
ÊܪJu�^�À>2 t�W��o � �W��o��>W�H�6J�L�6N�2��- �y�y.�>; u.�>su	�^�����D����Ȏ��+Y�>st������+6[�΋����@@�>su���������6o��� �>su������À>2 t+��W�� ��W�� �� ��� ��� Ë>W�L�6N�>; t�΋��AQS�VP�8��3ɋ.��8�>2 t�
�o � �
�o�� 렋6o�>a� �.]�6[�6Y��>; u�>su������� +��щk�.m3�Y�>; u�>st�������}�����
k+� ~
���+�Y�Y�}K�ًـ>; u�>	 u	�>s~u�&6k�������,6k��;>� r+>� ����6k�����
m+� ~)m~e�6m�c�y2�.�>s#t.8.;u.8.	t�����sP� ���X��u��&���& ���> �.�>; u.;>� r.+>� ��uڌȎ���P�ǀ� |��@|��`}��  XÁ�  X��P��H��X��P��.�@�� |��@|��`}��  XÁ�  X��P��H���3��28t��t38;t�	��������>s#u�Y�6[�J�6a�>; t� � �>s#u�Y�6[�(�6a�>; t� �%�b �>2 t�W��o � �W��o��>W�L�6N�����y�y.�>; u.�>su	�>�����$����Ȏ��� �>s~t��>2 t�J�o �	 �H�o��>o�]�� �ӡ�@@�>; u�>su������+���� �y�6a.�>s#tB.�>; t��.��������������u��5.�>su	� ����$�~ �;�r+�����o �r���vP� ���X��Ȏ�ø�+��]�>o�[�y�~8>�GGBu�3ۋY��y����+ڎy�6a��� �+�����y��P���Ȏ�ä�������Q.�����Q.���������Y�3�>2 tD�H�L;�}��>su+�= ����+�= } �Y�J�N+�}�؋J�6_��;�~�H$��Y�J�[3�����[ �]�Y�6[� �6aÀ>; t��.� �I�ޖ�>st�������>s~u�x�"2������ˊ���.� �>s#u�c ��t�d�����6� �&� �����6� ���3���9iu&>N�cË6� �>� �(�6� �>� ��6� �>� ������6� �>� ����;�|��;�~��À>�  t;� |;� ;� |;� �� ���À>9 t�R<`s���â�)��)�c)��)�g �� �W��o �y��
8"3��� �� �i�x�	�2��#u>� ��c�&f3��� ��@������ �� �� ��� ��� ��
U%���&u5� ��c�&f3��� �ءJ�Ɏ٣� �� ��� ����� �W��u��آs� ��c�&f3���.8&;tS��J�6c�ώ߉65�� �� �?�>; t�[�2�� �=P v	������� �� � ��   ��
8%��� ���&�&��sP�>; t��   ��s>��s5��s�>5t  � �g� �>; t�� � �� � ��&� �&�&�>; t�&>��g ��tB�>; u[��~t��
t���@t��tuG�����)��)�c)��)�&� �&� �� ��g  ���$t�>8 t�o�� ��� <t����	up�&� �&� �� `��d�f�� �����
&�g8&;t�y�&>��&� �&� �x�� �3��W��o���@�x�� �� ��>; t��@s
��w���r����d�f3��� ��8;u�� P ��t}�y ���u�i��	8;u(�.�/��
q"��
t%�3�>�W�>�o ?��t5�(r� �x�>; u$� �� �� �3E�WP�o��g �U�>; u�� ��� �g  �>j
qt9�y ��	�>; u(�.�/��
q"��
t%�3��W��o���u�>; u�3em�Wpm�on�� ^�� ��tQ�>; u�g S�� � �� ��� ��[uU�&2�>; u��.�/�y��
8"��
8%�� � �g  �>; u�� ��3��W��o���� �� ��0u:� �� ��� ^�� ��� 	�� 3��g�� ���Z�� �� ��� ���r� �>5�ut�>	 um�>5tf����"t��u�d��f�i ��d��!t��u=�d�f�g � �� ��� \�� ��� Z �� 	�� ���� �� �>5u/�>t(�02�U�� ��� ]��@����� ��2�������� �� H�>x t$��� �� H�� 3�8t��� 8&t��� �8&;t��� ��� �Fô� ���� ���� � ��� ��� ��� �2�8	t�8;u�
��=w��Ȏ�2�H������������� � �� ��]	�Ļ��ċ߹	 � ��Ļ0���>; u$�3� ��ڸ������ � B���J�Ĉ�Ɏٴ�)� � ��� �Z7p7�7�7)8G8�8_9�9�9�9�9�9�9�9�9�4
5
5
5
5
5
5
5
5
5
5
5
5
5
5
5
5
5
5
5�$4a4 �4[4 �R4�4	 �=4z4 �#4`4 ��4�4 ��4�4 ��4�4                                                                                                                                    O�4  �4 *** This is copyright 1984 Microsoft ***3��ء$0.�&�4����t<0u����t
��<0t���EÀ>7 t�SQR���� � �#4�t�`4���� � ��4�t��4� ��3ۜ����� � B�� � J��4�t��[4C��ٱ	�Ί��� � B�� � J��R4�t���4C��ٱ�4�� � ��<r ��t���� � B�� � ��=4�t��z4C�͋ٱ�4�� � ������ � B�� � J��$4�t��a4C��ZY[�P��$<	t<t�X��6�&�4��`t.��@��t;��@��t3��@��t*��@��t"��@��t��@��w	��r���2�������QW���>7 t,SR��3��4ڴ��
�t
��3��4�V� ��^Z[�\V��3�43����e����،Ȏ����4�< ���G�<+�������	�Z4��N�	��4��N���33���4��4@��4��4^3���� ���3������4�_Y�����r���wD�VP��% �����Ȏ����3X^π�w&.��4
�u.8&7uV�Ύފ�2��������3��4^�.�.�4��.��4P�~�X�3������3�� s�ÊËË�� ���3Ƅ�3���3s$2�� ���u�P�4��� � X���� � �����È��4��3��S�W�����33������s��_�W���ƅ�3���3���3���ێÎ�3����Q��s���Y+��%���u�P�4��� � X���� � P���X���G@��_�3����W��&�5���3&�E�������_�WR��&�5Ƅ�3���3���3&�E��&�e�$���u�P�4��� � X���� � P���X�����Z_�WRQS�؎���33�8otW�o�O��w����s���+��Ŋ$���u<t+���u<t"���u�P�4��� � X���� � P���X���F@�ƃ����3|�8.�4tN�.�4�W��4��4�� � � `4�#4�� � � ���� � �4�� � �>7 u�̠�4��4�� � �ʠ�4��4�[YZ_�WQ����2튍�38.7t��u��HTtI���3��4���3���ێÎ���s������Y_Ì؎���4�U��F�؋v�F]��.��4U��F�v�؉F]� �?������  ?  ���0���   @ ` p x | ~ � | l F                       ��  �?�F��������x�Ȏ�à:����>�:�:����>�#:à:����>�:�:����>�!:�P� ���:�:�%:����ڨu���&:����0�B�؊����u �%:�� ���:�İ�B�u�:�&:������	�B�J��$@�ǀt��u��:��B�J����@t��&:��t���H�:�:@�	8>:u��������� H�� ��B�J2�t���@t����B�:�:�.�:��~2����� @�� 3��x�!:�#:�� �� �*:�?����B�J
�t��B�t�*:�XË,:�.:�R����Z���ú��7�B���������7 �8��9 �:?�*:�(:�0�@�&*:�@���3 �@�@�@�Ë���3�9Ft�9Fu�F�?�F#�t�= w݋F#�t�= wѺ���B��PJ2���B��PJ2���B��PJ���B��PJ����B��PJ�����ĸ�B��PJ���B��PJ��ָ�B�J��P���B�J��P� ����~�>(:2��������Բְ���������&�&��θ ��v�ĸ�^��t(�N�~����������O����G����O�G������u��-�N�~������������O����G&�=���Ǫ��G������uӋ^�ְ0���@���^K@���X�X��X�X��X�X�X�X�X�Ë��5��&:��u��t���^�N���P�3���@���(:#�}+�3�@���@���1���X�þ���9�&��Ȍώǿ�9��ī����6��6�9�*:P��9P����á:
 �:��
;�wL�: �:��;�w;�B�@+F+D�>x t����BB������JӋ�_I���r�l��}���d��} �:+F�:+DRP�����Ë6!:�>:��6#:�>:�>:v+6F>F�m�:��.� �>�:�:��.� �>�:��� �D�F������ �������������7�B�$���������������<Ù�>� �<:�o��:�.�:��~2�����"%:�>u$�@��>���>� �>:�<��:�.�:��~2�����"%:�B�݋�+S+U���8t:��>t8;t�8>t%R����� � P���� � B�� � $�� � JX��Z��F�����BB������JӋ�_I�E휹 9t�J�.D�>�J�H�.B�>�H�9u�>x t�>H�øo�� ��� <@r<Ew������� ���� ��� �� �$�sP������� � B���X���5�� � P�	��� � B�<� � JX�>u�>> t8������>sw	�>sv�~���� � B���J�İ����� � B�� � $���V�Ύ�^�>u�>> t���L�������ꡅ�؊�A���ã� =P v	������� �� �� �?�g�� �D���� � ������ � B��
Ȁ�2�B�ËF��� ��>i������ ú��2�P�H�J���x�#�y���+�#�y���+ۀ� w< r� �>? t:@u	:Au�z�@�AU�������� � B�� � PJ���� � B�� � PJ���� � B�� � PJ���� � B�� � PJ��� � B�� � P��� � J���� � B�� � P2��� � J���� � B�� � P2��� � J�ΰ�� � B�� � P*����ǲĆØ��  �ˀ��ۀ� ������>c�ǿ����+��4�O����+��X������ � B���J�Ĳ�X������ � B���J��X������� � B���J��X������ � B���J������� � BX�� � J���� � BX�� � J���� � BX�� � J���?�� � BX���]��>? t���E�? �H#�y+ɋJ��<�t��#�y+ۺ��尜������ � B���J��@����� � B���J��@����� � B���J��@����� � B���J�İ��� � B�� � ��� � J�X��PQ��  �ȋŰ����� � B���J��H���� � B���J��H���� � B���J��H���� � B���J����YX#�tdPP���"�t!�ŋŬ�����Ŝ��� � B���J��H�ņ���"�t#���$N���Ŝ��� � B���J��H���Ȋ���uߪ*����"�tFXHu�XÜ������ � B�� � PJ���� � B�� � P2��� � J���� � B�� � P2��� � J��� � B�� � P�� � J���� � P��� � B�� � P*��� � J��� � B�� � P*��� � J��� � B�� � P*��� � J��� � B�� � P$��� � J��� � B�� � P���� ���� �ΰ�� � BX�� � J��� � BX�� � J��� � BX�� � J��� � BX�� � J��� � BX�� � JX��X������ � B���J��X������ � B���J��X������� � B���J��X������ � B���J�ĝòĀ>sw�>sv������ �`���� ������ �`���U��ދ������ � B���J�Ĺ  ��������K��s�]ÌȎغ����� � ����� � B좉�J���� � B���J�İ�� � B좊� J���� � B���J�İ�� � B�� � ��$�Ü�����&����� � B���J�İ�&����� � B���J�İ�&����� � B���J�Ġ��þ�
�u8
�t43�������؋��2�� ��ؿI�Ȏ��&�E �ЪG���Ȏ��z��H�Ȏ���3������������      X        ����  �   )P1P>PRP)P)P)P_PlP)P)P|P�P�P)P�P)P�P�P)P)P�P)PQQQ �Ȏ���35�!���t��3ɺHT�¸ �3�ǁ�HTu;ל�3�t�ǁ�HTu;�u�+G�6)G�?G�� ��6 �t��ʎں ru���l��� o3����PHu�8� ��؀>���u&�&tG�Ȏ�2�8/Gu�82Gt�80Gt�1G�>�1G
�u#�<�t)�<�t$�>0G u�1G
�u��2u
�� �� ��t׀�
����ع �<�u��:�u�������
JJ�m
�! ���r
�t��uK�>tG tD���
��;�
 �8tGt)��
��� ��
����r�
�t����	u��
 ��� �p������v��h���j
�Ո.k
�
�>� t@��Q�
�\�?���� � ����JJ�� � �BB�� � JJ�� � :�t�>0G u�� � �B��'2��� � 2�
�����
�uP� ��؀>����Ȏ�Xu��� �����u���uA��uA�����j
�k
��m
< j
�k
�>����R�� ��G�/G
�t��t�����D  �&��� �� s8�G�/G
�t��t�����D  ��� �.� �� �.� ����� �� � r���S�=�A뙴��
�u�&�G�q<�t�t<�t<�w��j
�0�!<r���t����>��.U��ʎº ��v���X+��>���s�����V��ŋ���~ u� ��h
���-G�3�j
�5�!�z
�|
���j
�%�!� ��ؿ�?�����4�xV�9��t � ��ظOL9J�t9P�t9�t9L�u.�&6�Ȏ���>5u� ��� � 3���u� � ����Atn�5� ����ͫu�:��3��ۈ�u^�-GG3�8;u89u�-G�9��-GS?���؊&I�c�ˎ���5�!��4��4�%��6�!�� 03ɋ���t�5�Ȏ��@ �&� ��y�.�  ��и5�!�r
�t
�%�h�!�35�!�v
�x
���3%�!�>9 t���6��6�9�*:P��P����� �>� t��x�-G� �G�O�G ��b�0�!����� �O3��G��s.� �G�� t��
u�GX �G����� � P�m
����B��R��
�� � �
J�Z� � ��
 ��R��
�Z"�2�"�t,��R��
�Z"�"�t�܊݊����s��C����u�Ȋ���2����R��
�ZXR��
�Z�í�m
��j
��k
�>m
 u�Ëm
��� � �P��� � �JJ� � �P2�� � �J� � �P�`� � ���� � �JJ� � �P2�� � �� � ��� � �J� � �P�= s"�m
X���X���BB����X�BX�BBX��g���
�m
B�����j
,��ð����3��؊l� � �:lt���� � �:lu��Ȏ؝��� � �J�� � ��Jθ 3��<u!��t��u�7�>= u� �>9 u�` ��B t%���
�u7&�Gt0�,:� �.:���0:�� u�H��2��B�$�<u	�9�-GS?Ë,:�.:����,:�0:���ø o���7Vu
�;�-GGø �3����KOu�5á� ���拴GWRV��	�!^Z��	�!�2�</tM<
t<u�2�.�>>G t8.83Gu2��@.8/Gt@.80Gt@.81Gt@.82Gt@��t��u@.84G����� 멠5G���6G"7G"8G<�t2������ �� �� �vƊ9G
�x2����2�8?Gt��>R t	�;G�.�3�<G
�x�.�3�6G"7G"8G<�t)� �3��86Gt�6G87Gt�7G88Gt�8G��3�9G
�x2�� �3�� �" �3�Ύư@�&� �y��. � �3�:G
�t2��- �3�Q�<
t<uNY�.�>G%� �؀�A��w���@G.�'Y���.�3G����� u�.�0G���� t�= w�.�/G
�t����.�8G.�� ���� .�6G.�� �� t�= w�.�1G���� .�� .��  �.�R� u��.�;G�� 
�t��.�<G.�Q�u��v��n �t�= w�.�:G��.�$.�"�U��Q u�= ~�.�9G�@��q .�7G.�� �o��c .�7G.�� �$�.�5G��� u�.�=���� u�.�2G���QR3ɋ���Ǹ
 ����s���u��؀�0r��	v�N��
�ZYù�������u�2 =d v�d �Q2���O ��<Ft+��<Nt+��<Dt��<St*����<Et��<Pt��<It2���N�Ċ�Y���� <Lt����
 <Fu�������<ar, �.�� .�� PSQRWVU�Ȏ��� ��
�>m
��F������ �>�wP���X������P������P2������������$��>� t�Ā�$$��
�2���t@��t��"� 
Ȉ� 3҈� �6@�>B�Ĩ t(�u�� �6� �>� �� ��� �6� �>� �� �t(�u�� �6� �>� �� ��� �6� �>� �� Y[�>� t�����.�� .�� PSQRWVU�Ȏ���>m
��FF�ְ��� � ���� � $��ְ��� � ���� � ��������
Ř�؋ְ��� � ���� � $��ְ��� � ���� � ����������
ŘP��3��� � �� ���Ћ6@�>B��������"���"� 
ц� 8� t&w�� �6� �>� �� ��� �6� �>� �� ���"���"� 
��� 8� t&w�� �6� �>� �� ��� �6� �>� �� Y.�� .�� PSQRWVU�Ȏ���m
�� � ������ � �����t�q
 �%�@u�>q
t�>q
t ����q
����q
� R��
�Z��� ���6@�>B3҈� �б��"���"� 
ц� 8� t&w�� �6� �>� �� ��� �6� �>� �� ��������"���"� 
ц� 8� t&w�� �6� �>� �� ��� �6� �>� �� ����������$��p
������o
��$?o
��
p
��Ƞo
����q
 ���� ��.�� .�� PSQ��·.�� �.�� s��u��t{���.�� �.�� s��uc��t_���.�� �.�� s��uE��tA��ˎûC&�� �&�� s��u"��t�ݸ ·&�� �&�� s��u��u��Y[X.�� .�� ø·.�� �.�� s��u���t���·.�� �.�� s���u���t���.�� .�� U��PSQRVW�Ȏ؋F�^
�N��2��
��4 � t�͉�2��t�ω�3҈� �Ћ6@�>B�"���"� 
ц� 8� t&w�� �6� �>� �� ��� �6� �>� �� �"���"� 
��� 8� t&w�� �6� �>� �� ��� �6� �>� �� ���_^ZY[X].�� .�� �.�� �.�z
.�>� u.�� �.�� PSQRWVU�Ȏ�������� �YW{W�W�W�WX%XGXiXbu�XPY�Z�\!_�ackdYf�gi�jl,o^p�r�u�X{Y)[]\_�a,c�dyf�g�i	kdlMo�p2sFv�X�Yd[Y]�_�aLc�d�f$h�i;k�l~o�p�s�v�X�Y�[�]�_
b�ce�fVh�i_k.m�oNq�s+w�XZ�[�]:`(b�cLe�f�hjk�m�o�qt�w�X@Z\^r`Vb�c�e"g�hCj�k�m�o�qKtxYpZK\Y^�`�b�c�eJg�hnj�k%n�or�t�x$Y�Z�\�^�`�bd�epg!i�j�k�n"phr�ty9Y�Z�\�^Ha�bCd.f�gVi�jl�nFp�r#uInvalid parameter
$Param�tre invalide
$Ongeldige parameter
$Ung�ltiger Parameter
$Ogiltig parameter
$Virheellinen parametri
$Par�metro no v�lido
$Par�metro inv�lido
$Parametro non valido
$Driver not installed -- Internal Error 1
$Gestionnaire non install� -- erreur interne 1
$Stuurprogramma niet ge�nstalleerd -- Interne fout 1
$Treiber nicht installiert -- Interner Fehler 1
$Drivrutinen ej installerad -- Internt fel 1
$Ohjainta ei ole asennettu -- sis�inen virhe 1
$Controlador no instalado - Error interno 1
$Controlador nao instalado - Erro interno 1
$Driver non installato - Errore interno 1
$Driver not installed -- Microsoft Mouse not found
$Gestionnaire non install� -- Microsoft Mouse introuvable
$Stuurprogramma niet ge�nstalleerd -- Microsoft Muis niet gevonden
$Treiber nicht installiert -- Microsoft Mouse nicht gefunden
$Drivrutinen ej installerad -- Musen kunde ej hittas
$Ohjainta ei ole asennettu -- hiirt� ei l�ydy
$Controlador no instalado -- El Mouse no se encuentra
$Controlador nao instalado -- Mouse nao encontrado
$Driver non installato - Mouse non trovato
$Driver not installed -- interrupt jumper missing
$Gestionnaire non install� -- cavalier
d'interruption introuvable
$Stuurprogramma niet ge�nstalleerd -- Onderbrekingsspringer niet
aanwezig
$Treiber nicht installiert -- Interrupt-Jumper
nicht gefunden
$Drivrutinen ej installerad -- avbrottsbygel finns inte
$Ohjainta ei ole asennettu -- keskeytyksen kytkin puuttuu
$Controlador no instalado -- El puente de interrupci�n no se encuentra 
$Controlador nao instalado -- jumper de interrup�ao nao encontrado
$Driver non installato - ponticello di interrupt mancante
$Driver not installed -- multiple interrupt jumpers found
$Gestionnaire non install� -- plusieurs cavaliers
d'interruption pr�sents
$Stuurprogramma niet ge�nstalleerd -- Meerdere
onderbrekingsspringers gevonden
$Treiber nicht installiert -- Mehrere Interrupt-Jumper gefunden
$Drivrutinen ej installerad -- multipla avbrottsbyglar
$Ohjainta ei ole asennettu -- liian monta keskeytyksen kytkint�
$Controlador no instalado -- Encontrados varios puentes de interrupci�n
$Controlador nao instalado -- m�ltiplos jumpers de interrup�ao encontrados
$Driver non installato - esiste pi� di un ponticello di interrupt
$MSX Mouse driver installed
$Le gestionnaire MSX Mouse est install�
$Microsoft MSX Mouse stuurprogramma wordt ge�nstalleerd
$Maustreiber MSX installiert
$Drivrutinen installeras Microsoft MSX MOUSE
$Asennetaan Microsoft MSX MOUSE laiteohjain
$Controlador MSX del Mouse instalado
$Instalando controlador da/do Microsoft MSX Mouse
$Installazione di Microsoft MSX Mouse Driver in corso
$Mouse driver installed
$Installation du gestionnaire 
$Microsoft Mouse stuurprogramma wordt ge�nstalleerd
$Maustreiber installiert
$Installerar drivrutiner f�r Microsoft MOUSE
$Asennetaan Microsoft MOUSE laiteohjain
$Controlador del Mouse instalado
$Instalando controlador da/do Microsoft Mouse
$Driver del Microsoft Mouse installato
$Switch values passed to existing Mouse driver
$Param�tres transmis au gestionnaire existant de la souris
$Schakelwaarden doorgegeven naar bestaand stuurprogramma
$Parameterwerte an vorhandenen Maustreiber weitergeleitet
$Parameterv�rden flyttade till existerande drivrutin f�r musen
$Kytkinasetukset siirretty olemassaolevaan ohjaimeen
$Par�metros transferidos al controlador en uso
$Defini�oes passadas para o controlador existente do Mouse
$Parametri trasferiti al driver esistente
$Existing Mouse driver enabled
$Le gestionnaire existant de la souris est activ�
$Bestaand stuurprogramma geactiveerd
$Vorhandener Maustreiber aktiviert
$Existerande drivrutin f�r musen aktiverad
$Olemassaoleva ohjain otetaan k�ytt��n
$El controlador en uso est� activado
$Controlador existente do Mouse ativado
$Driver esistente attivato
$Existing Mouse driver removed from memory
$Le gestionnaire existant de la souris est supprim� de la m�moire
$Bestaand stuurprogramma uit geheugen verwijderd
$Vorhandener Maustreiber ist aus dem Speicher entfernt worden
$Existerande drivrutin avl�gsnad fr�n minnet
$Olemassaoleva ohjain poistettu muistista
$El controlador en uso fu� retirado de la memoria
$Controlador existente do Mouse retirado da mem�ria
$Driver esistente rimosso dalla memoria
$Existing Mouse driver disabled
$Le gestionnaire existant de la souris est d�sactiv�
$Bestaand stuurprogramma inactief
$Vorhandener Maustreiber deaktiviert
$Existerande drivrutin inaktiverad
$Olemassaoleva ohjain poistetaan k�yt�st�
$El controlador del Mouse en uso est� desactivado
$Controlador existente do Mouse desativado
$Driver esistente disattivato
$Mouse Driver not installed
$Le gestionnaire de la souris n'est pas install�
$Stuurprogramma niet ge�nstalleerd
$Maustreiber nicht installiert
$Drivrutinen ej installerad
$Ohjainta ei ole asennettu
$Controlador del Mouse no instalado
$Controlador do Mouse nao instalado
$Driver non installato
$Mouse driver installed, cannot change port (/i, /z, /c, and /b invalid)
$Le gestionnaire de la souris est install�, impossible de changer de
port (/i, /z, /c et /b invalides)
$Stuurprogramma ge�nstalleerd, verandering van poort niet mogelijk
(/i, /z, /c en /b ongeldig)
$Maustreiber installiert, Anschlu� kann nicht gewechselt werden
(/i, /z, /c und /b ung�ltig)
$Drivrutinen installerad, kan inte byta port
(/i, /z, /c och /b ogiltiga)
$Ohjain asennettu, porttia ei voi vaihtaa
(virheellinen /i, /z, /c ja /b)
$Controlador del Mouse instalado,
no se puede cambiar el puerto (/i, /z, /c y /b no v�lidos)
$Controlador do Mouse instalado, nao � poss�vel mudar porta
(/i, /z, /c e /b inv�lidos)
$Driver installato, impossibile cambiare porta
(/i, /z, /c e /b non valide)
$Mouse driver already installed
$Le gestionnaire de la souris est d�j� install�
$Stuurprogramma al ge�nstalleerd
$Maustreiber ist schon installiert
$Drivrutinen redan installerad
$Ohjain on jo asennettu
$Controlador del Mouse ya instalado
$Controlador do Mouse j� instalado
$Driver gi� installato
$Unable to disable Mouse driver -- Control Panel is active
$Impossible de d�sactiver le gestionnaire de la souris --
le panneau de configuration est actif
$Niet mogelijk stuurprogramma uit te schakelen -- Controlepaneel is
geactiveerd
$Maustreiber kann nicht deaktiviert werden -- Steuerungsfeld ist aktiv
$Kan inte inaktivera drivrutinen -- Kontrollpanelen �r aktiv
$Ohjainta ei voi poistaa k�yt�st� -- ohjaintaulu on aktiivinen
$No se puede desactivar el controlador del Mouse-- El Panel de control est� activo
$Imposs�vel desativar controlador do Mouse -- painel de controle ativado
$Impossibile disattivare driver -- Pannello di controllo in
funzione
$Unable to disable Mouse driver -- Mouse Menu is active
$Impossible de d�sactiver le gestionnaire de la souris --
le menu souris est actif
$Niet mogelijk stuurprogramma uit te schakelen -- Muismenu is geactiveerd
$Maustreiber kann nicht deaktiviert werden -- Mausmen� ist aktiv
$Kan inte inaktivera drivrutinen -- Musmenyn �r aktiv
$Ohjainta ei voi poistaa k�yt�st� -- hiirivalikko on aktiivinen
$No se puede desactivar el controlador del Mouse-- Un Men� del Mouse est� activo
$Imposs�vel desativar controlador do Mouse -- Menu do Mouse ativado
$Impossibile disattivare driver -- Menu del Mouse in funzione
$Microsoft (R) Mouse Driver Version 7.04
Copyright (C) Microsoft Corp. 1983-1990.  All rights reserved.
$Microsoft (R) Gestionnaire de la souris.  Version 7.04
Copyright (C) Microsoft Corp. 1983-1990.  Tous droits r�serv�s.
$Microsoft (R) Mouse Stuurprogramma Versie 7.04
Copyright (C) Microsoft Corp. 1983-1990.  Alle rechten voorbehouden.
$Microsoft (R) Mouse Treiber-Version 7.04
Copyright (C) 1983-1990 Microsoft Corp.  Alle Rechte vorbehalten.
$Microsoft (R) Mouse drivrutin version 7.04
(C) Copyright Microsoft Corporation 1983-1990. Alla r�ttigheter reserverade.
$Microsoft (R) Mouse ohjainversio 7.04
(C) Copyright Microsoft Corporation 1983-1990. Kaikki oikeudet pid�tet��n.
$Controlador del Microsoft (R) Mouse Versi�n 7.04
Copyright Microsoft Corporation 1983-1990.  Todos los derechos reservados. 
$Microsoft (R) Unidade de Dispositivo Do Mouse Versao 7.04
Copyright (C) Microsoft Corp. 1983-1990.  Todos direitos reservados.
$Driver di Microsoft (R) Mouse Versione 7.04
Copyright (C) Microsoft Corp. 1983-1990.  Tutti i diritti sono riservati.
$Slow            Moderate        Fast            Unaccelerated   Faible          Moyenne         Maximale        Nulle           Laag            Gemiddeld       Hoog            Zonder          Niedrige        Mittlere        Hohe            Ohne            L�ngsam         Normal          Snabb           Oaccelererad    Hidas           Kohtuullinen    Nopea           Kiihdytt�m�t�n  Lento           Moderado        R�pido          No Acelerado    Devagar         Moderado        R�pido          Desacelerado    Lento           Medio           Veloce          Non accelerato                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             MZVQ W     ��    �rP`      �   ��L  �L  XM  �M  �M  �M  �M  N  N  )N  >N  �N  �N  �N  �N   O  O  }O  �O  �O  �O  Q  4Q  �Q  �Q  �Q  �R  �R  �S  HT  cT  �T  �T  U  'U  7U  @U  KU  RU  vU  �U  �U  �U  �U  V  zV  �V  EX  �X  �X  �X  "Y  HY  �i�����`�����_	��	��	��	��	��	�
�
�.
��
����������)�D�Y�m  m  �  ߊ  �  B�  ]�                                                                                                                                        ���� �lw12345678    OAK ATAPI IDE CD-ROM    ���c����������������E���2�������� T_ju��H����                                                                                                                                                                                                                             .�+ .�- �PSQRVWU�.� < t��.�+ �G�.�� �/ �G<v<�r,o<v�D�����t.�$�.�� 
�u��  ��N�u���Jr�!�!S.�� ��.���eu.��ft.Ǉf [����[���Kr��������D�T�|t�| t	�������O��Kr�����P�D�T�|t�| t	����������.��� .��� ����DT.;�H|.;�H|���� .��� .��� �Kr	.ƇT�L.ƇT 3�.��� .��� .��� .��� �53����������rs6�r1�1.��� .��� .;�� wr.;�� w.ƇT��Ks.ƇT ��3�.��� .��� .��� .��� .ƇT �Ը��c.��T��u������.��� .��� .��� .��� �@���c ��&�G8�v�����.�� .�$�� ��޸ ��l&�  &�M��W�sK_s�Z&�= t	&�=t�>�]&�E&�U���aK���K�W��K_r	&�&�U몸��� &�= t�0	&�=t3�&�E���Lr
&�&�U�{�3�&�&�U����L&��<�u"������3�.��� .��� .��� .��� .ƇT �r�<�����Mr�.���Nr�#���kNr���&�U&��&�MS&�]��[PSQRW��v� ��N_ZY[r$X��v���� ����� s	P�� ��X����3Y�7�wOr���,�OrDuN.��T�tK����&�����.��� .��� �:&�E&�U.��� .��� �%&�E&�U�k�.ƇT ���� .ƇT 3�&�&�E&�E&�E&�E���Qs�9�Or'P.�.� ����3�.��� .��� .��� .��� X���� &�<w�Or������o�Or�� ����b&�&�U&�u&�}��Or����I�Pr����?�Pr���5�Pr���+.�� �Pr���.�� � Pr������� �� .�+ �G.�  �v�]_^ZY[X�3��x s��[��3��| t@�|t��[���D�T�|tS.�� .��s�t.���t[�[�� VW��O_^s��[�� �L�\� �S.�� .ƇT [��VOË�.�� .��T�t�P�OXr.�� .ƇT ��u��[�9�SQ�؊�����	w������w	�	 �2�Y[��������
�����Q��2�����Ȋ���������Ћ�Y�S�؊±<��ǀ� �K ��2�Ã� -� �� [�Q� �� ����K���Y�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    ������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                        ������������������������������������������������                                                ffff                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                wwww                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        	5:   3     #6/    B}�d2��!:Sl���)[t��K                                                                                                                                                                                                                                                                                          � ����  s�.��H.��H���ʊ��.�>�H��t����P`  r�.�>nhuK.�Vh<t
<t<ts�9.�>`h(t*.�>`h)t"�'.�>`hu.��Hu�.�hc �-7�Q7u�.�>�H���u3��u��P`  � s� ��t� ��u� ���t� �� ���.��HtG� �P`  r>�!S��P`  [r,.�hc �6��6u�S.�� ��.Ǉ|e  [��  .�>�H��� �S.�� .���h [t�Ú�  s��  ��ʊ�д�t����P`  rø  ��Ú�  s���ʊ�д�P`  r���
��u���Ú�  s�v.��L �6O��.�T��.�D�ǋ��׸.���.�D���Ȏ�.������޴3ɚP`  ��r%.�W ��	r%<t<t.�Wu�
�P`  ����u��u����������Ú�  s�$�
�P`  .�W s����	r<u.�Wu������Ú�  s�
�"�P`  rø�����r�����t����.���
�u����<u�� �<u� ��3��.��.����.��;.��#�.��k.��S�.���.����Ú�  �&���.�d.�>b�z��Ӌ�C�P`  s&� �.�d.�>b��� �G�Ú�  �3�SQ�*.���h t�� ��� �P`  Y[s�� .���h u�e.��<pu�� <qu��.��� �u����� �u�������u���.��� �u������.��t���.�u���k.��<pu�� .��<qu��.��� �u����.��� �u�������u���.��� �u������.�t���.�u���Ʉ��3���.�>nhu.�Vh<u.�>`h(u����r�W���Ў����k s���_Ë�V�F��������  r"�.��[.Ƈ[ 
�u!��P`  s,.��[t� .Ƈ��.Ƈs��ñ�.Ƈ��.Ƈs�.Ƈ[ ����.�a ���/.�>nhu".�Vh<t<t�.�>`h(u�4.�>`hu�*���Ì�.�d.�>b��P`  r��.:��u�2.Ƈ���Ȏ���3ɻ��ʀ� t��$����  s뵴�P`  s�.�d.�>b.�� .���.�>a t�c3ɾ��ʀ� t��$�����D����ʀ� t��$���$�D����T��d��D����h t裴����踴.��H.��H��.�a���3�&�G���ʀ� t��$���Ȋ8�r@�D8�w9I��� ����T�d�DS.�� ���h [t�<�&�&�U�D���&�E�ø��Ú�  s�#.�U@�ӌȎؾYS�Ȏ��޴	�P`  [s����.�Ut�D<�tڱ��P� $<t3�X&�G�D��&�G�D&�G�T	�d
�D�t.���h t観�Ćª�«� ��T�d�D�t.���h t胳�Ćª�«����P��.�d.�>bX�����I�ʋЋ�.��L;�u
.��L;�u�.��L  .��L  ��QR���.��L�� .��LZY.��Lش&�P`  s�R�` ��ȋ�VW.�L.�>�L��@r�  .�>�L_^�s������.�d��.�>b�θ` ��ȾI����ø��Ú�  s��ӌȎؾf�Ȏ��޴�P`  s���ÊD��u���ÊD&�G�k�8���rK<tC��rB<u
.ƇT2��2�*<u
.ƇT2��"<u
.ƇT2��<u
.ƇT2��2�����Ú�  ����.�>�u�Ӹ�P`  r(�r#.�>� t���r��P`  ��.Ƈ��.Ƈs���Ú�  ���<t���P`  ��Ú�  s�)� �P`  ��P`  r�.�>`h)uS.�� .Ƈs�[�ø�Ú�  s�T.��.��;.���.��#��.��S.��k��.���.���.��.��;�
�t$
�t$.����Ӵ�P`  ����Ú�  r	�Ӵ�P`  ���������WS��  s�.�W
 .�Wu���FS�Ȏ�� 	3ɻY�P`  ��[r�.�E��������$<u�.�E
�u����� .�U.�e.�E[_��&r<u����SWV.��.��.����  s�n.�� .��s�uN.��H��㻻،Ȏ���P`  s���.�� .Ƈs �D�d.Ƈ� 8�t.Ƈ�R�	Zs�� .�� .���t� �� ��㾿��T�d�D���h t���<Kr,K�Ā�<r��<��.��.�&�.��.��.���� w��wr]<rY.:��wRr.:��wIr.:��w@<sK��,.��.��.�&�.��.�<Kr,K�Ā�<r��<��^_[.�����.��.��.��^_[�.�>nhu..�>`h(t.�>`hu.��Ht.�hc �,�,u�.�� ����.�� �� ��㾿��T�d�D���h t��<K|,K�Ā�<|��<���讋ʋ�.���O� ��P`  r5�O�<�u�<Cu�<Du�<0u�<0u�<1u�À��� �� �� ����Ú�  s�S���Ȏ���P`  r.��[�[�QS� � �*.�� .���h t����P`  rQ.��.�� .�&.���h t.�&.���h t�Ā���u.�� [Y��.�� .�&��t.���[Y�Q��  r>� � �*S.�� .���h [t�S���P`  [r�.�&���qt��pt� Y��Y��WQSPR���K�? 2��� I��� ��ZX[Y_ú? +ъ؈�WQP���K�? ��GI��G��XY_�WV.�0L  � ����ȌȎ؎��I.��K Q�� Q�Ȏ؎�� �VK�nK�Y.�2L.�.L��.�,L  �� .�,L��tQ�Ȏ؎�� �nK�VK�Y.�.L  �l.�,L��u	.�.L��t.�2Lu�.�0LW.�d.�>b�VK� ���r�tP+���X�Ȍ� ����.�d.�>b_..�KYIt�;��  .+0L^_�Q� �I��K�VK�2�.��L؁�@r��@݊$?&�G��.��L����@r�  .��LY�WVQS.��K .��K .��K .��K �VK� �������%�"�
�F2��.��K�VK� ��������
�F2��.��K�VK� ��������
�F2��.��K�VK� �$F�2���.�&�K.��K?u%.��K?u.��K?u.��K?u��.�,L ��.��K.��K.��K.��K.��K.��K.��K.��K� �3L.��L  .��K.2�K$?.��K.��K.2�K$?.��K.��K.2�K$?.��K.�>�K.�6�K�S��.�>�K.�6�K�D2��?�� u.�>�K u���ȈG.��K�G.��L�I.��K�.��K.��K����.��K.��K������.��K.��K.2�K$?.��K.��K.2�K$?.��K.��K.2�K$?.��K.�>�K.�6�K���.�>�K.�6�K�2��?�� u.�>�K u���ȈG.��K�G.��L�~It�_�.��K.��K.��K.��K.��K.��K.��K.��K� �3L.��L  .��K.2�K.��K.��K.2�K.��K.��K.2�K.��K.�>�K.�6�K���.�>�K.�6�K�
2��?�� u5���ȈG.�>�K.�6�K��.��K.2�K�������.��K2G.��LI.��K�.��K.��K��.��K.��K���.��K.��K.2�K.��K.��K.2�K.��K.��K.2�K.��K.�>�K.�6�K�l��.�>�K.�6�K�]2��?�� u5���ȈG.�>�K.�6�K�?.��K.2�K�d�����,.��K2G.��LIt�N�.�>�Lv�I�.�>�L u�>��3L�VK.��L2��G�G$?0 ���VK� �$F�2���.�&�K.��K?t���[Y^_�VQS.��K .��K �VK� ������� 
�F2��.��K�VK� �$F�2���.�&�K.��K?u.��K?t*.�.L �!.��K?t�� ��w�*�2��ؾVK.��K0 [Y^�W��K2�.��K��?�	.��K��?�)*�s��?_�$?��@t4$?�$?��s 4�$�$?�PSQ��?��?�߰ �ؘ��"��Թ �߰ �ؘ������"�2���Y[X�PV$?2�� ��K: t�����?*��K2��܊ ��^X�� �,0����������t��,0
Ī�� ������s�Ë� .Ƈ� .Ƈ��.�.���<Kr,K.���.�����S�
2������������[èu�u�u�u� �
������      ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            �                                                                          """"""""""""""""""""""""""""""""""""""""""""""""333333333333333333333333333333333333333333333333DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUffffffffffffffffffffffffffffffffffffffffffffffffwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwf3f3f3f3f3f3f3f3f3f3f3f3f3f3f3f3f3f3f3f3f3f3f3f3w3w3w3w3w3w3w3w3w3w3w3w3w3w3w3w3w3w3w3w3w3w3w3w3                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    � @p �� h
                                               	
pqrstuvw                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 �n�l|u�l�l�l�p�lvjwUxqx�x�l�l�x�xy�l�lUy�z�l�lXw�lo�l�lF{�uFwW{M|Nx)}t}�}o~���%��USQRWV��+�@ �ػ� �'��h ��h�.��g  �nh �oh �� �ph� �� �㋗�d��u��d��<f�>�g t�>�huB�hc� ���t	�$�<t����h ��g���>�k2���%2���P��X�.��h �^_ZY[]˴� �l�  ���l�  ����
��� ������ ���拔�c�P�[ X��$�<`u$�>nhu�>`h(t�>`h)uƇ[Ƈ��Ƈs��Ĩu��u�$�<u�n�< t�<0t�<Pt�<�t�<�t�<@t��z�S�� ���� �ph� ���g  �ph�th��g �E��s� �Th�ks� ���c�<t!S�뀿�h [t���d�tc�j���c�<tX�_���d�t�T��,d�B�������g��鋗lc�m��g9�gw��s�*S�뀿�h [t���d�t����c�<t�	���d�t[��nh��g+�g�ȃ� t�� �[Ë� �㋗�d�t�������g� �� ��� ��.��<f������g���c� ��B���hc ���u��hc� ��tB���d��<f�d�u"$�<Pt< t<uۋ�\d�<�t�	J�<u�������d��<f4�� ��^c0	�\c �Kb���g  ��g  ��g  ��g  �Vc�Xc3Ҹ0	�&Xc��g��g3��Zc�ph��qh S�� ���h t
�ph��qh [��g�rh��g�sh��g�th��g�uh�Xc�vh �&wh�xh�yh��zh ���g� �� ��3Ҹ0	�>Xc~	S� ��[��&Xc��ઊ�<f�����s� �Ks�%����c�<t&S�뀿�h [t���d�u� �b����c�<tv�V����d�t�����\d��J���g��g Q�Yt`��g��g;�gu;�gt�yrM눀>Hbu���r9S�뀿�h [t���d�t������c�<t������d�t��t�e��;���j��Q��l��^c �\c �Kb �Ib �Hb �>Vc u�k�>Mc u�a���f u���f t���Hb�H�@ ���{  u�	�``� �D  �����fc �Vc�`c�bc�``�(s�fc��s�\c�Vc��bc�Vc�s
<Ut�����S�M�� u	�Mc  ���]f�f�Gs t�ЋG+D���Tf�fG3�f���G�D������[�>fc t�Vc)bct�^c�&Vc���	�p����L ��`c�Vc��`�}
 u��r[�Mc��gf�Ef�Mc�\g���<fu&�F��Ib���.fPfQfW�``� �D  �����Vc�Xc3Ҹ �>Kb t�0	�&Xc��`��`f�    f�    �>Pc�Rc�f��fǨt	f_fYfX�� f��`�``� Qf��`f�f�>�`   r,f3�+ȉL�� uf�   f�`f)�`��Y��f_fYfX�Yf�>�` u���.�`s"t �С�`+D���Tf��`f�`3�f����`�D�L �f�    �ȱf��f``  �Mc��gf�Mc�\g���<fu&�F� � ��Ib�f_fYfX�>Ib u
�>Kb t�����g  ��g  ��g  ��g  ��h�Vc�Xc3Ҹ �>Kb t�0	�&Xc��g��g3��Zc�ph(��g�rh��g�sh��g�th��g�uh�Xc�&wh�xh�>Kb t�ph��yh��zh ���g��>Ib u� �� ���>Kb t3Ҹ0	�&Xc�3Ҹ �>Xc~	S� ��[��&Xc���.��<f�����es�!�>Ib u�.�Mc�\g���<fu&�F� � �Mc�,g�	� � �� ��s�����c�<t)S�뀿�h [t���d�u� ������c�<t���� ���d�t�~���\d��J���g��g Q�'Yu� ��g��g;�gu;�gt��s� �G��S��>Hbt(�>Ib t$�Mc�,g�$�� � ��@ ���{  t�^�f�rVS�뀿�h [t���d�t�E����c�<t�9����d�t%�����>Ib t�)�@ ���{  t��t���t���������ph+��g�rh��g�sh��g�th��g�uh��g  �bS�� ���h [t�E��
r5�r8���c�<t���hc� ��t���d���h�t��h �;�t������#��&
��h ��g ��h@���h ��g ��h ��g  �phC�qh��h�vh��g�&wh�xh��h�yh��g��g��>
s�� �>Pc�Rc��
s�� ���c�<t�����d�t����\d��J���� tA�g��鋗lc�ă���g��g t��gI�����g9�gtL�|
s� ���c�<t�����d�t�K���\d��J���� tA�g��鋗lc�����g9�gt��0
r7S�뀿�h [t���d�t�V����c�<t�J����d�t���t����������h��g ��h �"��h��g ��h@���h��g ��h@�phB�qh��h�rh��h�sh��g�&wh�xh��g��g�a
��s� �h�	s� ���c�<t�����d�t�V���\d��J���g��鋗lc�m��g9�gu��F	rUS�뀿�h [t���d�t�l����c�<t�`����d�t���>Pc�Rc�h��g�>�h t�h�����t��������h���h �phK��h�xh��g  �	���s����g �sh�6Pc�Rc�Ɏ�� �ɎٰG�ph�� ���h t� �sh���	����g  �H	�`�ph�qh �th ��g  �-	�E�ph�qh �th��g  �	�*�ph�qh �th��g  ���� �>�g u���>�gr����ph�th �>�gt
�ph�th��g  ���� ������phU�qh�rh �wh �xh��g ��g ��g ��g ��g ��g � h �h �h�h�h�h �h �h �h �	h �� � �� t
������� �
h���h� ��; t
���#��� �h��;�h���S���h ��k�h�������h ����h����g ���Ys�v��g���rp���c�< t�,􋗼d�t���\d��J���g�����lc�o�>�gr��r4S�뀿�h [t���d�t����c�<t��󋗼d�t�z�t�[��e��.��ph�th$��g$ �:�rl�>Pc�Rc�`rg���c�<t�󋗼d�t�2�\d��J���g��鋗lc�m��g9�gu��"r)���c�<t���d�t�J󋗼d�t���t���������ph ��g  �����g  �phZ��g�rh��g�wh��g�xh�&�g��g��g��s� �>Pc�Rc�s� ���c�<t#S�뀿�h [t���d�tm����c�<ta�򋗼d�t�U�\d��J���g��鋗lc�m�Nr\���d�t	���c�<t�S�뀿�h [t���d�t�b��c�<t�V򋗼d�t���t����g+�g�ȃ� t�� ��������g  �ph�th��g ��"s� �>Pc�Rc��s� ���c�<t#S�뀿�h [t���d�td����c�<tX��񋗼d�t�p���\d��J���g��鋗lc�m��g9�gw��`rJS�뀿�h [t���d�t���c�<t�z񋗼d�t��t����g+�g�ȃ� t�� �������trB���d�����r6���d�u� ��lc����!���c�u���\d�<�t�J�<t��u���t����g� �� ��� ����<f�����r/��r'���d�u�>Pc�Rc� ��鋗lc�m�h�(���'��U��ph%��g �2�s� �fh�Xs� ���c�<t�����d�t�'\d��J���g��鋗lc�m��g9�gu��rGS�뀿�h [t���d�t�=����c�<t�1����d�t���>Pc�Rc�fh� ��~�t����Vc�Xc3��Zc��g  ��g  3Ҹ` �&Xc��g��g�ph��qh �zhS�� ���h t�ph��qh �zh@[��g�rh��g�sh��g�th��g�uh�Xc�vh �&wh�xh�yh ���g� �� ���` �&Xc��ઊ�<f�����{s� �"s��틗�c�<t#S�뀿�h [t���d�tx�<�c�<tl�0�d�t��틗\d��J���g��g Q�zYtV��g��g;�gu;�gt�KrC��r9S�뀿�h [t���d�t���c�<t���d�t�h�t�I�����N��5��P����g�Jb����g�� �� ����<f����s����$�:r���d�u����Jbt������������i r4�r7S�뀿�h [t���d�t�9�c�<t�-�d�t���t������&�g��g�.�g��g�6�g��g�Pc�Rc�>Vc�6TcË� ���rM���lf u�� r<���c�<u7���d�t.��- r#���c�<u���d쨀t����ph� ��lc�o��2������� r)�hc .�>~h�t�hc� �c�t���d�$�<t���Ë��d���S��hc �4S� �hc6 �(S�� � ���hc� &�� ��&���eu�hc���)t0��hu�1<u��@ �ػ� ��t�'�����h �� [���� [�Ë��d;��duQ�� ��Y�hc .�>~h�t�hc� ���t���d쨀u������hc .�>~h�t�hc� �y�t���d$�<@u��������g� �� ����g��ઊ�<f��������g���c� ��B���PSQR�䡊�� �!�� �㋗lc�> ��#��!��� ��ZY[X�PSQR�䡊�� �!.�� ��.��lc� ��!��� ��ZY[X�V� ��h.;t����^��.�L^��VSQR.�� ��.��lc� ��h.;t������.�D�ZY[^���`� �E  �``�E�E  �ȉE�< ����Krf�E�@�����`�Vc�Xc3Ҹ �>Kb t�0	�&Xc��E  �Pc�u"�E�E  �Rc�E�E �E  �  ����KðU��À>Kb u	�>bc r�Ã>bcr������`����  �K��P��� � 䠨t
� �� � � X���P�!.�|h� �.�}hX���P.�|h�!� .�}h�X��SQ��g��g��g��g3�3�3���gXc��g��Kr0��K��g��g����Ks��g��<r��<��g��g����<s��g��g�&�g��gY[À�ds	��<s<Ks ��S�Pc�Rc�؀?ds�<s�Ks�ds
�<s�K�Ȏ��[ÜPS�@ �ۻl ��_.�jc.hcs.�jc[X��PS�@ �ػl ��_.;jcr	.;hcr3�[Xù S�
2�����������Ī��[�Pcs�Pcs�Rc �Ë>Pc�Rc���r�tP+��
 X�Ȍ� �����lc��>Hb t��f�m��m��SRVP�w�2�6�h�P�5�!��g��gX�%�`��!�@ �ػ� �'X^Z[�PS�>�ht��g���$��h�)�<r� �� � � � R.�� ���d�Z[X��VRP���2�6�h�%.��g.��g�!XZ^��RVPS���2�6�h�P�5�!��g��gX�%���![X^Z�PS�>�ht��g���"��h��<r� �� � � R.�� ���d�Z[X��VRP�n�2�6�h�%��g��g�!XZ^�RVPS�I�2�6�h�P�5�!��g��gX�%����![X^Z�PS�>�ht��g���"��h��<r� �� � � R.�� ���d�Z[X��VRP���2�6�h�%��g��g�!XZ^�RVPS��2�6�h�P�5�!��g��gX�%���![X^Z�PS�>�ht��g���"��h�z�<r� �� � � R.�� ���d�Z[X��VRP�R�2�6�h�%��g��g�!XZ^�   .�hc	 �����u���ph��xh �yh(��g( �l���g  ���s�u�>Pc�Rc��rp���c�<t���c�<tJ�拗�d�t�S勗\d��J���g��鋗lc�m��g9�gw��C�r)���c�<t���d�t�k拗�d�t��t����������ph��qh �th&�� ��&��Le�&wh�xh��g  �����PSQRV&�� ��&�� &��Le t&���eA��J&��Le t���;&���eA&��|e�����ھ &���eA&��'t.Ƈ[.Ƈ��.Ƈs�C����^ZY[X�SQ�� �ph� ���g  �ph��xh �yh(��g( ����s�o�'�<�rg���c�<t���c�<tG�S���d�t�H��\d��J���g��鋗lc�m��g9�gw����r"���c�<t���d�t����d�t����Y[�PSQR&�� ��&���et�6�< �8�sPSQRW���_ZY[X��&�'����&�'�`t	�������ZY[X�SQS&�� &���h [t� �*��� � �P`  s�
&�$�<�t�Y[�PSQRWV&�� P��2��X2��I��}&�� K��&Ǉ�e � � ��S&�� K��&ǇLe  &��|e&���e&Ǉ�e [P&��lc&��<f&�� ��&��<fX&��lcB&���cB&���c��&��,dB&��\dB&���dB&���d&��lc��&���dB&��e&�� &��Le&��|e&���e&Ǉ�e @�^_ZY[X�PSQR�< S�'�(�P`  [sS�'�(�P`  [r&�'���V�&�'�`t	�g������ZY[X�PSQR&�� ��&���et�A� &��Le&;�|eu�1�)�P`  s.�Vh<u
.�>`h:u�	�)�P`  s��e�r��u���ZY[X�SV� �I�r&�� ��&��Le����&��'��u�p�� ^[�PSR�� �㋇Le��,d�|e��\d��� ����X[Z�                fPSRf�Ӌ���@f�� � � ��f�f�׋�� ����f���af��뀿�fu#f�Ӌ���Df�� � � ��f�f�ߋ��f���af�f�Ӌ���f�� � � ��f�f�ۋ�� �〿�f tf���f���f��f3�f�Z[fX�fPRf�Ӌ���@f�� � � ��f�׋f�f�Ӌ���f�� � � ��f�ۋf��f3�f�ZfX�         � �
          

This driver is provided by Oak Technology, Inc..
OTI-91X ATAPI CD-ROM device driver, Rev D91XV352
(C)Copyright Oak Technology Inc. 1987-1997
   Device Name        :    
  Number of drives   :  

 
  Invalid /p switch  :  
  No drives found, aborting installation
 
  Transfer Mode      :  Programmed I/O  PCI Bus Master DMA 
  Firmware version   :    Port=    IRQ=  
  Drive   12345678 AB                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��p�p���h�h�                   S�  ��.�� �w�<t
<
t</t����.�� � <bu�l<su�<dt<pu�O<vu�<qu�뼃�� �
 �< t<t<
t<	t���NQ�� t� ���X� +ȃ� u� .���}��|:t1F� <iu%� <ou.���<0r<4w$.�.��J�N�F����^s�<�< u�Rrw�ж �Ir���
���< u�8��<,uY.���*s< t��I���sN���	��w8u
.��.�>�u�2��h� &;t�����&�G�ȸ ��&�G� ����.���2��< u����<,u�<0u���<1u ��.����.����.��.��.���N�F� <mt�.�� .���<0r<2w$.� .��놊��� ��su	.���s��s�.���g�.���^�[.���
 ��&�.�FG������ �.�>� u����� �� .������ ��rf.��&�Mcf.��f&�Ӌ.�>�t .�>�u �s	�  ���;.�>� u"����%� �?&�>Mc t&�>�f t�O� .��&� �  ��s����� �n 3��  &�& ���G�W�G �G rF.�>� u)����� �@ &� ��
rRQ3��±
����r YZ���k .�>�t�.�>� u������ � �PR.�G"�t��!��ZXì<0r <:r<Ar<Gr<ar<gs,W��,7��,0���Ã�r��w������RP��
r��7���0��!XZ�.�>�u��VPSQR.�� .�� .�� .�� .�� .�� .�� .�� .�� �6�&��   � .�>�u� &�~h��&�� �㬊ଋЬ&��<f&��lcB&���cB&���c��&��,dB&��\dB&���dB&���d&��lc��&���dB&��e&ǇLe  &Ǉ|e  &Ǉ�e  &Ǉ�e  �3� �P`  s��QR&���d&��<f�� � � JJ��� � � �U�� � � � � � �<U� � � ���ZYt���#�P`  s��r��S���$�P`  [s�.�����t�����t�x$`< u&Ƈlf&�>Mc u�� �s�� .�>�t.�>� tV.�1 uO.�1 tD.�>u.�&��g�.�O t'&��g.�O t&��g�'�P`  r	&Ƈ�f���h.�� .�� .�� �*.�>� t
.� .���#.�>�u.�K�r*�.��.�M�r.�� &��g�'�P`  r��&Ƈ�f ��P`  ��P`  S����P`  [r&��<u�
�P`  ���  s�FS�'�(�P`  [s�6&�&'��&�,. ����  &���f t�*�R�&���f t�.�B�
.��&�� �� ��It.�>�t�z�.�>� u�������&�~h ZY[X^�S�z��P`  ��[r1&�=u+&�}Nu$&�}	Eu&�}
Cu&�} 3sS&�� &Ƈ�h[����`2�.���  Q������7����}��:��!�|�&��lc��&����d��ր�����������T��ր��L��������hQ2�&�&9�lct����Y&�D<
r��!�,
������CY�a�&��e���u.���"��wu.������u.���.���&��e���u.�>� uV�#�  .���I��wu.�>� u;�Å  .���.���u.�>� u �Q�  .���.�>� u�߆  .���&��e���u.�>� uV���  .�� �I��wu.�>� u;�.�  .�� �.���u.�>� u ���  .�� �.�>� u�J�  .�� ÜPS�@ �ۻl ��_.��.�s.��[X��PS�@ �ػl ��_.;�r	.;�r3�[X�&��e���u.&Ƈ�f&Ƈ,g &Ƈ\g&Ƈ�g.�� &��<ft.���2��wu.&Ƈ�f&Ƈ,g&Ƈ\g
&Ƈ�g.��&��<ft.������&��e���u.�� ���wu.�����èu
�u�u��.����.����.�� ��PSQ2��I���:���Y[X�PSQ2��I��&Ƈ�f��Y[X�fPSQ2��I��f&���a��f&���a��Y[fX�&���d�t
&���dnt�&���d��&���d� � � �8�t�&���d&���d�          � ���       fRSQP����r-.��.�����t�) .�>��u.��t�1.�>��uXY[fZ��XY[fZ��RfP��f.��f�� � � ��f�� � � f=t|f=�ttf=��0tlf=��ptf=��qu&��g�T.�.�.�>��u��8WSQ2۹@ �>Mbf.���ú�f�� � � ��f�� � � f&�������Y[_��f3�f�fXZ�.�>��u�f.��f.�����f�� � � �����t���.��f.�����f�� � � �����t���.��f.��� ��f�� � � ��f���f.���C�RP���� ��=t4=�t$=��t�� 2Ҁ��u��2��XZÀ��=0t����=t�ր��=u�.�>��uв .������t���.������t���.���"�f�������f.����  �  �  ��  ��  ��    �  �  �  ��  ��  ��   	      @   �   �   �  �  �  ��  ��  ��    �  �  �  ��  ��  ��                   @   fPQVf.�����@f�� � � ��f�6�.�>�u�6@.�>� tf%��  ���f%  ��.�>� t��3�.�������f.�kr/fPS�6(.�>�u�6p�.�>� t��f.���f&���a[fXS��f&���a[^YfX��  �  �  �  0�  0�  0�  0�    �  �  �  �  0�  0�  0�  0�fPRVf.�����@f�� � � ��f�.�>� tf%��  �f%  ���6+.�>� t�� &��<ft��.�>u#.�>r)��.�>t��.�>t�����&�>�gt��f.�` rOfPS�6(.�>u.�>v��.�>t�����&�>�gt��.�>� t��f.���f&���a[fXS��f&���a[^ZfX�&�>�gu&&��<ft.�>� uf @  �f   @&Ƈ�f����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          MZ�C V     ��      �E      ;   "2  Q2  �2  �2  �2  33  Q3  a3  t3  �3  �3  �3  4  "4  K4  V4  �4  �4  5  .5  e6  6  �6  ,7  77  &8  I8  19  �9  �9  (:  ?:  [:  r:  �:  �:  �:  �:  �:  ;  $;  /;  @;  j;  �;  �;  �=  �=  �=  >  m>  �>  �IY�!	=	�	B
N
U
`
r
w
�
�
>Yt������P  �P  �m  �n  �n  ;o  Vo                                                                                                                                            ���� �� � 12345678    OAK ATAPI IDE CD-ROM    eee�eee=eeee�GVee=eQ��=ee�ee49>Vp�����;F��)3                                                                             .�+ .�- �PSQRVWU�.� < t��.�+ �G�.�� �/ �G<v<�r,o<v�D�����t.�$�.�� 
�u��  �N�u���0r�!�!S.�� ��.��Ju.��<Jt.Ǉ<J [����[��1r��������D�T�|t�| t	�������O�1r�����P�D�T�|t�| t	����������.��� .��� ����DT.;Z.|.;X.|���� .��� .��� �s1r	.Ƈ� �L.Ƈ�  3�.��� .��� .��� .��� �53����������rs6�r1�1.��� .��� .;�� wr.;�� w.Ƈ� �1s.Ƈ�  ��3�.��� .��� .��� .��� .Ƈ�  �Ը��c.��� ��u������.��� .��� .��� .��� �@���c ��&�G8�v�����.�� .�$�� ��޸ ��l&�  &�M��W�N1_s�Z&�= t	&�=t�>�]&�E&�U���<1���1�W��1_r	&�&�U몸��� &�= t�0	&�=t3�&�E���2r
&�&�U�{�3�&�&�U����2&��<�u"������3�.��� .��� .��� .��� .Ƈ�  �r�<������2r�.����3r�#���F4r���&�U&��&�MS&�]��[PSQRW��v� ��4_ZY[r$X��v���� ����� s	P�� ��X����3Y�7�R5r���,�5rDuN.��� �tK����&�����.��� .��� �:&�E&�U.��� .��� �%&�E&�U�k�.Ƈ�  ���� .Ƈ�  3�&�&�E&�E&�E&�E����6s�9�b5r'P.�.� ����3�.��� .��� .��� .��� X���� &�<w�v5r������o�5r�� ����b&�&�U&�u&�}�5r����I��5r����?��5r���5��5r���+.�� ��5r���.�� ��5r������� �� .�+ �G.�  �v�]_^ZY[X�3��x s��[��3��| t@�|t��[���D�T�|tS.�� .����t.���t[�[�� VW��5_^s��[�� �L�\� �S.�� .Ƈ�  [��15Ë�.�� .��� �t�P�5Xr.�� .Ƈ�  ��u��[�9�SQ�؊�����	w������w	�	 �2�Y[��������
�����Q��2�����Ȋ���������Ћ�Y�S�؊±<��ǀ� �K ��2�Ã� -� �� [�Q� �� ����K���Y�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    ��������������������������������                                                                                                                                                                                                                                                ��������������������������������                                ffff                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                wwww                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        	5:   3     #6/    B}�d2��!:Sl���)[t��K                                                                                                                                                                                                                                                                                          � ���o  s�� .�W..�S.���ʊ��.�>T.��t�����E  r�.�>&LuK.�L<t
<t<ts�9.�>L(t*.�>L)t"�'.�>Lu.�W.u�.�xH �q5�5u�.�>T.���u3��u���E  � s� ��t� ��u� ���t� �� ���.�S.t2� ��E  r)�!S�m��E  [r.�xH �5�%5u�.�>T.�*�� �S.�� .��cL [t�Úo  s��  ��ʊ�д�t�����E  rø  ��Úo  s���ʊ�д��E  r���
��u���Úo  s�v.�2 �6���.�T��.�D�ǋ����.���.�D���Ȏ�.������޴3ɚ�E  ��r%.�� ��	r%<t<t.��u�
��E  ����u��u����������Úo  s�$�
��E  .�� s����	r<u.��u������Úo  s�
�"��E  rø�����r�����t����.���
�u����<u�� �<u� ��3��.���.����.���.����.��.����.��#.���Úo  �&���.��.�>�����Ӌ�C��E  s&� �.��.�>���� �G�Úo  �3�SQ�*.��cL t�� �O� ��E  Y[s�� .��cL u�e.�Q<pu�� <qu��.�[�� �u����� �u�������u���.�\�� �u������.�[�t���.�]u���k.�Q<pu�� .�Q<qu��.�\�� �u����.�[�� �u�������u���.�^�� �u������.�]t���.�]u���Ʉ��3���.�>&Lu.�L<u.�>L(u����r�W���Ў����k s���_Ë�V�F�+Ѓ����o  r"�.���.Ƈ� 
�u!���E  s,.���t� .Ƈ��.Ƈ���ñ�.Ƈ��.Ƈ��.Ƈ� ����.�� ���/.�>&Lu".�L<t<t�.�>L(u�4.�>Lu�*���Ì�.��.�>����E  r��.:��u�2.Ƈ���Ȏ���3ɻ3�ʀ� t��$���o  s뵴��E  s�.��.�>�.�� .���.�>� t�c3ɾ5�ʀ� t��$�����D��3�ʀ� t��$���$�D����T��d��D���cL t��Ϋ������.�X..�Z.��.�����3�&�G�5�ʀ� t��$���Ȋ8�r@�D8�w9I��� ����T�d�DS.�� ��cL [t�a�&�&�U�D���&�E�ø��Úo  s�#.��@�ӌȎؾ�S�Ȏ��޴	��E  [s����.��t�D<�tڱ��P� $<t3�X&�G�D��&�G�D&�G�T	�d
�D�t.��cL t��͆Ćª�«� ��T�d�D�t.��cL t�͆Ćª�«����P��.��.�>�X�����v.�ʋЋ�.�2;�u
.�2;�u�.�2  .�2  ��QR���.�2�� .�2ZY.�2ش&��E  s�R�` ��ȋ�VW.2.�>2��@r�  .�>2_^�s������.����.�>��θ` ��Ⱦv.����ø��Úo  s��ӌȎؾ��Ȏ��޴��E  s���ÊD��u���ÊD&�G���8���rK<tC��rB<u
.Ƈ� 2��2�*<u
.Ƈ� 2��"<u
.Ƈ� 2��<u
.Ƈ� 2��2�����Úo  ����.�>Nu�Ӹ��E  r(�r#.�>M t���r���E  ��.Ƈ��.Ƈ����Úo  ���<t����E  ��Úo  s�)� ��E  ���E  r�.�>L)uS.�� .Ƈ��[�ø�Úo  s�T.���.���.���.�����.���.����.��.��#.���.����
�t$
�t$.����Ӵ��E  ����Úo  r	�Ӵ��E  ���������WS�o  s�.��
 .��u���FS�Ȏ�� 	3ɻ���E  ��[r�.�E��������$<u�.�E
�u����� .�U.�e.�E[_��&r<u����SWV.�.�.��o  s�n.�� .����uN.�V.����،Ȏ����E  s���.�� .Ƈ� �D�d.Ƈ� 8�t.Ƈ�R�	Zs�� .�� .���t� �� ������T�d�D��cL t�ʱ�<Kr,K�Ā�<r��<��.�.�&.�.�.��� w��wr]<rY.:�wRr.:�)wIr.:�9w@<sK��,.�.�.�&.�.<Kr,K�Ā�<r��<��^_[.����.�.�.�^_[�.�>&Lu..�>L(t.�>Lu.�V.t.�xH ��*�+u�.�� ����.� �� ������T�d�D��cL t��<K|,K�Ā�<|��<���ɋʋ�.���� ���E  r5���<�u�<Cu�<Du�<0u�<0u�<1u�À��� �� �� ����Úo  s�S�I�Ȏ����E  r.�J[�[�QS� � �*.�� .��cL t��O��E  rQ.�N.�� .�&].��cL t.�&[.��cL t�Ā���u.�N [Y��.�M .�&]��t.�M�[Y�Q�o  r>� � �*S.�� .��cL [t�S�O��E  [r�.�&Q��qt��pt� Y��Y��WQSPR��1�? 2��� I��� ��ZX[Y_ú? +ъ؈�WQP��L1�? ��GI��G��XY_�WV.��1  � ����ȌȎ؎��v..��0 Q�� Q�Ȏ؎�� ��0��0�Y.��1.��1��.��1  �� .��1��tQ�Ȏ؎�� ��0��0�Y.��1  �l.��1��u	.��1��t.��1u�.��1W.��.�>���0� ���r�tP+���X�Ȍ� ����.��.�>�_..�0YIt�;��  .+�1^_�Q� �v.��0��0�2�.�2؁�@r��@݊$?&�G��.�2����@r�  .�2Y�WVQS.�1 .�1 .�1 .�1 ��0� �������%�"�
�F2��.�1��0� ��������
�F2��.�1��0� ��������
�F2��.�1��0� �$F�2���.�&1.�1?u%.�1?u.�1?u.�1?u��.��1 ��.�1.�1.�1.�	1.�1.�
1.�1.�1� ��1.�2  .�1.2	1$?.�1.�	1.2
1$?.�1.�
1.21$?.�1.�>1.�61�S��.�>1.�61�D2��?�� u.�>1 u���ȈG.�1�G.�2�I.�	1�.�	1.�
1����.�
1.�1������.�1.�1.2	1$?.�1.�	1.2
1$?.�1.�
1.21$?.�1.�>1.�61���.�>1.�61�2��?�� u.�>1 u���ȈG.�1�G.�2�~It�_�.�1.�1.�1.�	1.�1.�
1.�1.�1� ��1.�2  .�1.2	1.�1.�	1.2
1.�1.�
1.21.�1.�>1.�61���.�>1.�61�
2��?�� u5���ȈG.�>1.�61��.�1.21�������.�12G.�2I.�	1�.�	1.�
1��.�
1.�1���.�1.�1.2	1.�1.�	1.2
1.�1.�
1.21.�1.�>1.�61�l��.�>1.�61�]2��?�� u5���ȈG.�>1.�61�?.�1.21�d�����,.�12G.�2It�N�.�>2v�I�.�>2 u�>���1��0.�22��G�G$?0 ����0� �$F�2���.�&1.�1?t���[Y^_�VQS.�1 .�1 ��0� ������� 
�F2��.�1��0� �$F�2���.�&1.�1?u.�1?t*.��1 �!.�1?t�� ��w�*�2��ؾ�0.�10 [Y^�W�12�.�1��?�	.�1��?�)*�s��?_�$?��@t4$?�$?��s 4�$�$?�PSQ��?��?�߰ �ؘ��"��Թ �߰ �ؘ������"�2���Y[X�PV$?2�� �L1: t�����?*�L12��܊ ��^X�� �,0����������t��,0
Ī�� ������s�Ë� .Ƈ .Ƈ)�..��9<Kr,K.��9.��)��S�
2������������[èu�u�u�u� �
������           �U
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            �                                                          """"""""""""""""""""""""""""""""33333333333333333333333333333333DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUffffffffffffffffffffffffffffffffwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwf3f3f3f3f3f3f3f3f3f3f3f3f3f3f3f3w3w3w3w3w3w3w3w3w3w3w3w3w3w3w3w3                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            � @p �� h
                                       	
pqrstuvw                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 >R�P,Y�P�P�PeT�P�Y[\!\o\�P�P�\�\�\�P�P]g^�P�P[�P�R�P�P�^�Y�Z_�_�[�`$atabuc0k�k�USQRWV���@ �ػ� �'�[L �\L�"��K  �&L �'L �� �(L� �� �㋗|I��u�<I��\J�>�K t�>�LuB�xH� ��t	�$�<t����L ��K���>�O2���%2���P�X�.�\L �^_ZY[]˴� �em  ���em  ����
��� ������ ���拔�H�P�[ X��$�<`u$�>&Lu�>L(t�>L)uƇ�Ƈ��Ƈ���Ĩu��u�$�<u�n�< t�<0t�<Pt�<�t�<�t�<@t��z�S�� ���� �(L� ���K  �(L�,L��K �9�s� �L�_s� ���H�<t!S�뀿cL [t��\I�tc�j���H�<tX�_��\I�t�T���H�B�������K��鋗|H�m��K9�Kw���s�*S�뀿cL [t��\I�t����H�<t�	��\I�t[��&L��K+�K�ȃ� t�� �[Ë� �㋗\I�t�������K� �� ��� ��.��\J������K���H� ��B���xH ���u��xH� ��tB��<I��\J\I�u"$�<Pt< t<uۋ�I�<�t�	J�<u������<I��\J4�� ��nH0	�lH �[G���K  ��K  ��K  ��K  �fH�hH3Ҹ0	�&hH��K��K3��jH�(L��)L S�� ��cL t
�(L��)L [��K�*L��K�+L��K�,L��K�-L�hH�.L �&/L�0L�1L��2L ���K� �� ��3Ҹ0	�>hH~	S� ��[��&hH��ઊ�\J�����s� �?s�%����H�<t&S�뀿cL [t��\I�u� �b����H�<tv�V���\I�t�����I��J���K��K Q�Yt`��K��K;�Ku;�Kt�mrM눀>XGu�[�r9S�뀿cL [t��\I�t������H�<t�����\I�t��t�e��;���j��Q��l��nH �lH �[G �YG �XG �>fH u�k�>]H u�a���J u���J t�7�XG�H�@ ���{  u�	��E� �D  �����vH �fH�pH�rH��E�s�vH��s�lH�fH��rH�fH�s
<Ut�����S�M�� u	�]H  ���]f�f�Gs t�ЋG+D���Tf�fG3�f���G�D������[�>vH t�fH)rHt�nH�&fH�����p����L ��pH�fH�8F�}
 u��r[�]H�TKf�Ef�]H�4K���\Ju&�F��YG��.fPfQfW��E� �D  �����fH�hH3Ҹ �>[G t�0	�&hH�4F�6Ff�    f�    �>`H�bH�f��fǨt	f_fYfX�� f�0F��E� Qf�0Ff�f�>4F   r,f3�+ȉL�� uf�   f0Ff)4F��Y��f_fYfX�Yf�>4F u���.4Fs"t �С4F+D���Tf�0Ff4F3�f���4F�D�L �f�    �ȱf��f�E  �]H�TKf�]H�4K���\Ju&�F� � ��YG��f_fYfX�>YG u
�>[G t�����K  ��K  ��K  ��K  �`L�fH�hH3Ҹ �>[G t�0	�&hH��K��K3��jH�(L(��K�*L��K�+L��K�,L��K�-L�hH�&/L�0L�>[G t�(L��1L��2L ���K��>YG u� �� ���>[G t3Ҹ0	�&hH�3Ҹ �>hH~	S� ��[��&hH���.��\J�����Ys�!�>YG u�.�]H�4K���\Ju&�F� � �]H�K�	� � �� ��s�����H�<t)S�뀿cL [t��\I�u� ������H�<t���� ��\I�t�~���I��J���K��K Q�Yu� ��K��K;�Ku;�Kt��s� �G��G��>XGt(�>YG t$�]H�K�$�� � ��@ ���{  t�R��rVS�뀿cL [t��\I�t�E����H�<t�9���\I�t%�����>YG t�r�@ ���{  t��t���t���������(L+��K�*L��K�+L��K�,L��K�-L��K  �VS�� ��cL [t�E��
r5�ur8���H�<t���xH� ��t��\I���L�t��L �;�t������#��
�^L ��K �_L@��^L ��K �_L ��K  �(LC�)L�^L�.L��K�&/L�0L�_L�1L��K��K��2
s�� �>`H�bH��
s�� ���H�<t����\I�t����I��J���� tA�K��鋗|H�ă���K��K t��KI�����K9�KtL�p
s� ���H�<t����\I�t�K���I��J���� tA�K��鋗|H�����K9�Kt��$
r7S�뀿cL [t��\I�t�V����H�<t�J���\I�t���t���������]L��K �aL �"�]L��K �aL@��]L��K �aL@�(LB�)L�aL�*L�]L�+L��K�&/L�0L��K��K�U
��s� ��K�{	s� ���H�<t����\I�t�V���I��J���K��鋗|H�m��K9�Ku��:	rUS�뀿cL [t��\I�t�l����H�<t�`���\I�t���>`H�bH��K��K�>aL t��K�����t�������bL��bL �(LK�bL�0L��K  �	��s����K �+L�6`H�bH�Ɏ�� �ɎٰG�(L�� ��cL t� �+L��������K  �<	�T�(L�)L �,L ��K  �!	�9�(L�)L �,L��K  �	��(L�)L �,L��K  ���� �>�K u���>�Kr����(L�,L �>�Kt
�(L�,L��K  ���� ������(LU�)L�*L�/L �0L��K ��K ��K ��K ��K ��K ��K ��K ��K��K��K��K ��K ��K ��K ��K �� � ��� t
������� ��K�����K� ��� t
������� ��K�����K��������K ����K�������K ��#��K����K ���Ms�v��K���rp���H�< t�,�\I�t���I��J���K�����|H�o�>�Kr��r4S�뀿cL [t��\I�t��󋗼H�<t���\I�t�z�t�[��e��.��(L�,L$��K$ �.�rl�>`H�bH�Trg���H�<t��\I�t�2�I��J���K��鋗|H�m��K9�Ku��r)���H�<t��\I�t�J�\I�t���t���������(L ��K  ����K  �(LZ��K�*L��K�/L��K�0L�&�K��K��K�w��s� �>`H�bH�s� ���H�<t#S�뀿cL [t��\I�tm��򋗼H�<ta��\I�t�U�I��J���K��鋗|H�m�Br\��\I�t	���H�<t�S�뀿cL [t��\I�t�b򋗼H�<t�V�\I�t���t���K+�K�ȃ� t�� ��������K  �(L�,L��K ��s� �>`H�bH�s� ���H�<t#S�뀿cL [t��\I�td��񋗼H�<tX���\I�t�p���I��J���K��鋗|H�m��K9�Kw��TrJS�뀿cL [t��\I�t�񋗼H�<t�z�\I�t��t��K+�K�ȃ� t�� �������hrB��\I�����r6��\I�u� ��|H����!���H�u���I�<�t�J�<t��u���t����K� �� ��� ����\J�����r/��r'��\I�u�>`H�bH� ��鋗|H�m�\�(���'��U��(L%��K �&�s� �L�Ls� ���H�<t����\I�t�'I��J���K��鋗|H�m��K9�Ku��rGS�뀿cL [t��\I�t�=����H�<t�1���\I�t���>`H�bH�L� ��~�t����fH�hH3��jH3Ҹ` �&hH��K��K�(L��)L �2LS�� ��cL t�(L��)L �2L@[��K�*L��K�+L��K�,L��K�-L�hH�.L �&/L�0L�1L ���K� �� ���` �&hH��ઊ�\J�����{s� �"s��H�<t#S�뀿cL [t��\I�tx�H�H�<tl�<\I�t��틗I��J���K��K Q�zYtV��K��K;�Ku;�Kt�KrC��r9S�뀿cL [t��\I�t���H�<t��\I�t�t�t�U��+���Z��A��\����K�ZG���|K�� �� ����\J����s����$�:r��\I�u����ZGt�����������i r4�r7S�뀿cL [t��\I�t�E�H�<t�9\I�t���t�������&�K��K�.�K��K�6�K��K�`H�bH�>fH�6dHË� ���rM���|J u�� r<���H�<u7��\I�t.��- r#���H�<u��|I쨀t����(L� ��|H�o��2������� r)�xH .�>6L�t�xH� �c�t��|I�$�<t���Ë�\I���S��xH �4S� �xH6 �(S�� � ���xH� &�� ��&��Ju�xH���)t0�[Lu�1<u��@ �ػ� ��t�'����[L �� [���� [�Ë�|I;�\IuQ�� ��Y�xH .�>6L�t�xH� ���t��|I쨀u������xH .�>6L�t�xH� �y�t��|I$�<@u��������K� �� ����K��ઊ�\J��������K���H� ��B���PSQR�䡊�� �!�� �㋗|H�> ��#��!��� ��ZY[X�PSQR�䡊�� �!.�� ��.��|H� ��!��� ��ZY[X�V� �9L.;t����^��.�L^��VSQR.�� ��.��|H� �9L.;t������.�D�ZY[^��8F� �E  ��E�E�E  �ȉE�< ����Krf�E�@����HF�fH�hH3Ҹ �>[G t�0	�&hH��E  �`H�u"�E�E  �bH�E�E �E  �  ����KðU��À>[G u	�>rH r�Ã>rHr�����HF����  �K��P��� � 䠨t
� �� � � X���P�!.�4L� �.�5LX���P.�4L�!� .�5L�X��SQ��K��K��K��K3�3�3���KhH��K��Kr0��K��K��K����Ks��K��<r��<��K��K����<sK��K�&�K��KY[À�ds	��<s<Ks ��S�`H�bH�؀?ds�<s�Ks�ds
�<s�K�Ȏ��[ÜPS�@ �ۻl ��_.�zH.xHs.�zH[X��PS�@ �ػl ��_.;zHr	.;xHr3�[Xù S�
2�����������Ī��[�`Hs�`Hs�bH �Ë>`H�bH���r�tP+��
 X�Ȍ� �����|H��>XG t��f�m��m��SRVP�w�2�6sL�P�5�!�~K��KX�%�i�!�@ �ػ� �'X^Z[�PS�>\Lt�~K���$�[L�)�<r� �� � � � R.�� ��\I�Z[X��VRP���2�6sL�%.�~K.��K�!XZ^��RVPS���2�6sL�P�5�!��K��KX�%��i�![X^Z�PS�>\Lt��K���"�[L��<r� �� � � R.�� ��\I�Z[X��VRP�n�2�6sL�%��K��K�!XZ^�RVPS�I�2�6sL�P�5�!��K��KX�%�%j�![X^Z�PS�>\Lt��K���"�[L��<r� �� � � R.�� ��\I�Z[X��VRP���2�6sL�%��K��K�!XZ^�RVPS��2�6sL�P�5�!��K��KX�%��j�![X^Z�PS�>\Lt��K���"�[L�z�<r� �� � � R.�� ��\I�Z[X��VRP�R�2�6sL�%��K��K�!XZ^�               .�xH	 �����u���(L��0L �1L��K �`���K  ��K �Q����s�u�>`H�bH�u�rp���H�<t���H�<tJ�拗\I�t�J勗I��J���K��鋗|H�m��K9�Kw��.�r)���H�<t��\I�t�b拗\I�t��t���������(L��)L �,L&�� ��&���I�&/L�0L��K  ����PSQR&�� ��&�� &���I t&���IA��J&���I t���}&���IA&���I������&��t.Ƈ�.Ƈ��.Ƈ��C&��t.Ƈ�.Ƈ��.Ƈ��C&��t.Ƈ�.Ƈ��.Ƈ��C&��t.Ƈ�.Ƈ��.Ƈ��ZY[X�SQ�� �(L� ���K  �(L��0L �1L��K ���B�s�o����rg���H�<t���H�<tG�S��\I�t�H��I��J���K��鋗|H�m��K9�Kw���r"���H�<t��\I�t���\I�t����Y[�PSQR&�� ��&��Jt�6�( �8�sPSQRW��_ZY[X��&����j�&��`t	�r������ZY[X�SQS&�� &��cL [t� �*�O� � ��E  s�
&�]$�<�t�Y[�PSQRWV&�� P��2��X2��I��}&�� K��&ǇJ � � ��S&�� K��&Ǉ�I  &���I&���I&ǇJ [P&��|H&��\J&�� ��&��\JX&��|HB&���HB&���H��&���HB&��IB&��<IB&��\I&��|H��&��|IB&���I&�� &���I&���I&���I&ǇJ @�^_ZY[X�PSQR�< S��(��E  [sS��(��E  [r&�����&��`t	�������ZY[X�PSQR&�� ��&��Jt�A� &���I&;��Iu�1�)��E  s.�L<u
.�>L:u�	�)��E  s��e�r��u���ZY[X�SV� �I�r&�� ��&���I����&����u�p�� ^[�PSR�� �㋇�I���H��I��I��� ����X[Z�                fPSRf��o���@f�� � � ��f�f��o�� ����f���Ff��뀿�Ju#f��o���Df�� � � ��f�f��o��f��Gf�f��o���f�� � � ��f�f��o�� �〿�J tf���f���f��f3�f�Z[fX�fPRf��o���@f�� � � ��f��of�f��o���f�� � � ��f��of��f3�f�ZfX����z          

  CD-ROM Device Driver for IDE (Four Channels Supported)
  (C)Copyright Oak Technology Inc. 1993-1996
  Driver Version     : V340
  Device Name        :    
  Number of drives   :  

 
  Invalid /p switch  :  
  No drives found, aborting installation
 
  Transfer Mode      :  Programmed I/O  PCI Bus Master DMA 
  Firmware version   :    Port=    IRQ=  
  Drive   (Primary Channel)  (Secondary Channel)  (IDE Channel 3)  (IDE Channel 4) , Master , Slave  12345678 AB                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              ��p�p���h�h�                  S�  ��.�� �w�<t
<
t</t���.�� � <bu�d<su�<dt<pu�G<vu�{�Ã�� �
 �< t<t<
t<	t���NQ�� t� ���X� +ȃ� u� .��녃|:t1F� <iu%� <ou.���<0r<4w$.��.���R�N�N����s�D�< u�rw�ж ��r���
���< u����<,uY.����s< t��I����sN���	��w8u
.��.�>�u�2�9L� &;t�����&�G�ȸ ��&�G� ������.���2��< u�v��<,u�<0u���<1u ��.����.����.��.��.���N�F� <mt�.�� .���<0r<2w$.��.����.���{�[.���
 ��&�.�FG���� S��  �O��� � � �[���� � .����� �	rf.��&�]Hf.��f&��o.�>�t .�>�u �� s	�  ��3�����n �3&�>]H t&�>�J t�C�U .��&� �  �s����� �; 3��  &�& ���G�W�G �G r.��.�>�t�������� � �PR.�G"�t��!��ZXì<0r <:r<Ar<Gr<ar<gs,W��,7��,0���Ã�r��w������RP��
r��7���0��!XZ�.�>�u��VPSQR.�� .�� .�� .�� .�� .�� .�� .�� .�� �6�&��   � .�>�u� &�6L��&�� �㬊ଋЬ&��\J&��|HB&���HB&���H��&���HB&��IB&��<IB&��\I&��|H��&��|IB&���I&Ǉ�I  &Ǉ�I  &Ǉ�I  &ǇJ  �[� ��E  s��QR&��<I&��\J�� � � JJ��� � � �U�� � � � � � �<U� � � ���ZYt��-�#��E  s��r��S���$��E  [s�SQVW�Ȏ������� ���� ��%G�GFF��_^Y[.�����t�����t�M$`< u&Ƈ|J&�>]H u� �s� .�>�t.�>� t	.�� uF.�>�u.��&�|K�.� t'&�|K.� t&�|K�'��E  r	&Ƈ�J���F.�� .�� .�� �/.�>� t
.��.���	.��r.�� &�|K�'��E  r�����E  ���E  S�I���E  [r&�J<u�
��E  ��m  s�FS��(��E  [s�6&�&��&��. ���m  &���J t�Q�y�&���J t�U�i�
.��&�� �"��It.�>�t�y�.�>� u�������&�6L ZY[X^�S�����E  ��[r1&�=u+&�}Nu$&�}	Eu&�}
Cu&�} 3sS&�� &ƇcL[����`2�.���  Q������6����|��:��!�p�%��|H��&����c��ր�����������S��ր��K����y����9LQ2�&�&9�|Ht����Y&�D<
r���,
��������V���� ��� S�����[����CYI�� t�a�a�&���I���u.���"��wu.������u.���.���&���I���u.�>� uV��h  .���I��wu.�>� u;�gi  .���.���u.�>� u ��i  .���.�>� u��j  .���&���I���u.�>� uV�Ai  .�� �I��wu.�>� u;��i  .�� �.���u.�>� u �`j  .�� �.�>� u��j  .�� ÜPS�@ �ۻl ��_.��.�s.��[X��PS�@ �ػl ��_.;�r	.;�r3�[X�&���I���u.&Ƈ�J&ƇK &Ƈ4K&ƇTK.�� &��\Jt.���2��wu.&Ƈ�J&ƇK&Ƈ4K
&ƇTK.��&��\Jt.������&���I���u.�� ���wu.�����èu
�u�u��.����.����.�� ��PSQ2��I���:���Y[X�PSQ2��I��&Ƈ�J��Y[X�fPSQ2��If&���F��f&���F��Y[fX�&��|I�t
&��|Int�&��\I��&��|I� � � �8�t�&��\I&��|IÜ�|H&� =�t=pt=�t=ht�������������������\J&� <�t<�t�������������             � ���       fRSQP����r-.��.�����t�) .�>��u.��t�).�>��uXY[fZ��XY[fZ��RfP��f.��f�� � � ��f�� � � f=ttf=�tlf=��0tdf=��pu&�}K�T.�.�.�>��u��8WSQ2۹@ �>]Gf.���ú�f�� � � ��f�� � � f&�������Y[_��f3�f�fXZ�.�>��u�f.��f.�����f�� � � �����t���.��f.�����f�� � � �����t���.��f.��� ��f�� � � ��f���f.���C�RP���� ��=t4=�t$=��t�� 2Ҁ��u��2��XZÀ��=0t����=t�ր��=u�.�>��uв .������t���.������t���.���"�f�������f.����  �  �  ��  ��  ��    �  �  �  ��  ��  ��   	      @   �   �   fPQVf.�����@f�� � � ��f�6�.�>� tf%��  ���f%  ��.�>� t��3�.�������f.�gr#fPS�6�.�>� t��f.���f&��G[fXS��f&���F[^YfX��  �  �  �  0�  0�  0�  0�    �  �  �  �  0�  0�  0�  0�fPRV�3�f.�����@f�� � � ��f�.�>� tf%��  �f%  ���6�.�>� t�� &��\Jt��.�>�u#.�>�r)��.�>�t��.�>�t�����&�>|Kt��f.�d rOfPS�6.�>�u.�>�v��.�>�t�����&�>|Kt��.�>� t��f.���f&��G[fXS��f&���F[� �^ZfX�&�>}Ku&&��\Jt.�>� uf @  �f   @&Ƈ�J����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          �����W;�si��-D�%������ ��~��ر����S3�S�PKLITE Copr. 1992 PKWARE Inc. All Rights ReservedNot enough memory$� 	�a�!� ����OO����������FF� ��� �2�����;����<����A����c����d����e����f���r���Jt�s�3�3���Jt�����Jt��Ӆ�t��Jt��Ӏ�r��Ju�����.����
t:3ۃ�t&��Jt�r��Jt�����Jt�����Jt��Ӏ�s.��,���V��+��^눬Ȁ� <�u��3��Ju����Ӏ�r���Ju����Ӏ�r���Ju����Ӂ�� ���3�� S�؋ȋЋ����� 
      	          	
�  �-�Converted  MZ L @    �� d��B�,���  RJ%0;)�FQ\g�Rr}�J)��������E'V�$�%QR&+rJI��'I��)A*������-���	.����0$%%39�cEQ4�6�8RR��9E�;=>�CQ�}D�E�$GK%)LD�P��EQ�R���q�t w �Q  �Y R7 ����� ��w � Bi��ں�!� ,�	%�0НU�6 BZ,�o^�`�"M� Me7bB�n0ȜG�X2 G��B>�$7[�!�{�u�,	]�
Hu]�u]�u]�u]�u]�uM� ]�!"#��$y�ԥ%&X[�T'(u])*+p�k�H-�.u]$/01�n2c<��3n4u}$56ЭT�08�9:;��<� ���,9�
u�F0G
=u0I]�KLM�[N��O���P���Q0R��0S0T��0U0VW�<X<Y<Z��[C������] 
:($6MS DO  Version 6 (C)Cop (yright 1981- T94 MicrosofA�rp Lensed� at;ial - %"P!p&yթ &/Al�Mse2r�Lv5� �FMT.EXE �B	�K� �#/;G  S_kw�����%������f2	} � 
Oض	/VB?S��41:8B Pn�G	�T���NTELECT:5ACKUPA �UTOTES$�
�uFU]?QC8� T �
@P
! #~!��JA����)(����������� ���R
���J)@���N�	@	J)��� %+0m 160K%�B88,L320;3K-�K7igK<��0Kd�.2M��440K��!�EM28Ng�K��.M�B%o*?[  ]:<|>+=;,/\."()&-�^����j����R]�>o�]r f:\-�L�zn.? �.A:CONA�3PH�xx�(�F)<CFg�� �
̑@
��� 
�"��:\I0�O.SYS
MS�hNO NAM:E�	F�D�'�0 ���Ȏ�3ҎҼ |(
��` ����  �ri� r�.�>|t�h.�d}� N�Q�	*�� ��(V-3���.�6����ƴ<-^Y.� )6|t.�&e}@���űQ��.;T�|G���
Qu�g}��� P2�.�$tV�� 	�^����3�u� S�Yr3���&� M�H  G����}@���u� �	�þ`�� ����
Non-S pystem disk or�
errRe 
place and %ri�*ky �when�adycP& D9Boot fail�_u�,Inc io��'sr0msdn �w/��~ �� u�~�;uv@#��]�7��Q<�,5.0F�/Qb��g��	�GkU� 	JFAT12�3�� ���x 6ŀ7VS�>|^  ��E��|�M��G�����y�59|t  � |�|�&|H@||�� �P�R|�IK|� 
 $|� �H(���� �'� .� r�������}�X 
� �t��( }�_ �^��D( �X��GHH�@�|2���Z, ZY� PRQ�%:Q�XT YZXrH	� ���� K.|�$�4�3�p �
�t�)���;� �s�6�O|�R3�|
% U�M|���ô�@�
���
6�ʆ�hQ�6!�$M�p�s#�IOC[�����q��B�#�9S��6	�l'
�s���A:���H=FO�RMAT,�r�p ���=:`�@ @��(>��:S	>h�b� `	�ա�]��J]>@�WR>��$l��� �^Iv�
�;��Q��iW -�X:\CO {MMAND.h���uSPEC=�(@DRVACE.BIN�K7i=P߽����-S�wtack!-��  PSRW3Ɏ�3��.�  ��/���>�)m��S������%)�������״M�--	 ���
�M

$	  P�
 ��8mR����R
.A  (Q�P rY_Z[XG �����PV� c�!B��6�{�^X��D�3�P�����D��R �0=u�� �= s�����
�  �B� �� fSQUWR���6 (���t�u
& 0�Z�L�_����
Z�r]Y��DEA?����
5,5wo�YlY��2�6	�t;�tR Ir��� �u�&�-��$E� sUUM�H� 	GIu���WP (S���ٰ��� H+�K��[X_�3�-	SOA�@��Z(��UP=�Z X�X�B� P&�=u����� ��UQ����YsJa�ȩ;��* "]q�' � �PÀ���ƀu  ~�>� � ��W�> �&�= �t& :r�:Ew�GG�  �_Ï3ۓ��6����	v��7�
0RA�uB�t 9�u�|
,u�6P�A�"]�c �3�맨Re� 	!�%� &8%
`u
et:�u 
S�s�BI u�V���t3M�>f�u+�D0�A*��<0��6@�4��>fuBP 4IOO����W+�� (
�_Ys��Q�ʊH� tu#TQ�^�u�	�:3�TVgQ'(
m-�DSP�|�tnt��B� � �z`N  rY_]^�p
�Dr8$��c�%� (i��X��C��@�(0�����
�TC���VS3��� �h����ߠ@�%��tu���È-p=' i�w����&(�7���p�����t��� tlT ��Ȣ�r����  +u)RUQWP� �/ 	<�Xu	�ظ��T�s_�\��� ]Z�[^߹Z2 X����I�E(\G�Z��t=uP��
�l ��t&�M�	 Q.85u.��Ld-��@%&;�.�	� I���r�@�&}Q@�2�FG�� U��u`�: -CCƢ
C覭3�
 �$�D	:�v*����t
�|| ��u��E8Ls*B��ъ�$��S��7Aa�A;�u�B�Uu
�Y#�YEBC�
�t &d��u���U�x��#ˬ�>9�Z�r��p$��]60uxPAH �@�s�EP��c bGA�!�+�D]�TUX H"4 u$"Qp�u��C$p�v�u�	�T�u&&'
�*��+C�,��
,(&n[U*�*�O 	*@t)PR�82Th��ҨL�,���ZX�,��TA�ǈ	����BN��-R���( ��G��k�L��   � K k	 �(g� �� P  5 R  �o � � �   �Z [ �,{-  �.�/$0`1� �2��4 �5T6�7�8  j9C:z;�<���=%���orrect;~�v�@�
*%1 �W���"mpleted.	��B*byb�v�ab+ �XC�(zH,F_ma D��
CI
�Ji@bad)��?s�tal��1sp�T(#�)�(rbnew*�e( fD)Vri� :]U:Zu,X�%����!Rei�@<.Volu��m�ez(1��Jchar{*l�, ENTER3�n�e)? $�*�supp�B:�� T0�v�i��devid��pRdS»Lrom)�3r.1 Ey IOT�CTL�>l.PR<Npa�M�lock?. ?�!BwSt2FFg:.~!d$iry/��Can�f�� ASSIGN��3SUBST���V0U�0JR�FilesM!PM�tw��k@"$�a jj(�v�%\��DQ��|bX�0��-#Tod��,� th�r� /��O:mX�oif(sM[S��aM(I{ou� �^BL^n@,ad.)���
WARNING: _��)nta&�,eV�me�\Aa�<�r���Ywil��!troyos�	=<�n;�fӛ�
y|��]P?�1�O F(��ywa%(Y/N)?'9�dp��n��1MS-�ʧG?�] z`��[/V[:�]]4MQU`F:size
B | /��S
C]@LT@T:t$k�Ґ�:1�MM�1]�4@9@
z�388+  Ǧ m�pp��ifixq0�c5�,Q �Per� �jq��uick�RG)1)U
)n u!�nd��)�2F2��j77�of�loppy۟�t@(such��=��a@160,8dN32�7
1.244)2.88)�GuB�B >Al[�a�6l�$��|x�`������H:HS HC�}��%v��L.�� 2nuX8mber
#\!��lideycf>�N!?J;�77;1 � )�E[ngleSCb<a��M8�/4
85.25-<h�tK+�, P�high-TnYtyO��0N8.uNe,t��?1C 1T-X`!clusVC�����u�*EntljP"rko"P��."@#�	��	  H  a  �    �  �   7   O j � � �  �# �$  % 4& B' c( �B�P 2�jOHg�h�mina�G�Z��un]it�/��� Peʍa��T;Vt 0�-���Cus�A1UnL��k@	BOOT.�¸�Z ��N.�argetwQs�d�� C#�� [�A. �+��ID.����nsf{*�e*���nfM[ ��aI .�8�ati��H=4Ѹx �!#Y�"t�� tJ��SQi��N�n-%2�P b1�Hkeܥ��[�� �y�L�y~B�P��aT� *���� �%) � * � + � ,- � .
  / ?0 ]1 {2 �  3 �4 �5 �6   7 :8 w9 �: '  ; �< F 8G a  K uL �M �N Z  O hP vQ �R �  S T U $V @ �W ^X qY �%d�@G�.Wy��Qcm#a�"2^�A
�LL'ATA ON N (-REMOVABLEXISK)DRIVE$�WI+BL��UT!x#�qEa�o�Fhr!-w!�"�#�Dr��a���5unitVS	�)#����;�7� ��S� J[`�tw�$�Mx�@p���i5(/NA��)@TryoԵD�ZS���CAie
MrouUQgn�S �ScsT2�a\st����swY&<�4b!�O�UNz.�4�k- ��8zsLĲw�� ��d@
 <f]z��t#��o�T*�G;cQ�����7C�t���u��%8�#��xЊy/i�2u3�i&;�2���4�N,�ufb�~ci�ay`��lo-�lc
�-rQ�	��kԾEx��\�s݊ԟ7-�5�\h�e�tX�k�	[U5?�iF��c%1K X�M#�.%2v����y��ZR�Zg�sh���Vfy{���P�|�v�w�i��a�heck~x"p��u� =�-
p	s�=  ��8� f19'197  B G1j/��y �R B J�Too2�ny op� �KAc#Ec	�t �	�[:�BLK+T�tyExt=�aP5)и�J�(U� ����C�W; �"����N��RVW����͎����u�  �]�u�M�u�U	��8}
���_^Zi��ÛV� []|<>+=;" P@.�m�.�`�tbu:�f1��6J
;@�f�s�S&��B&:s�\�#(N6oSWU�wU  �n uC���r<�Z�t7�u�"lP�&AtN� 
0�<=u.�C����bŬC�NTWd ���$	st�6`�</t6"tGu 
T&�G2�.9�s
(.���CC�2`+� �i�	�J`(@��2�CSQS'��sAl�4��,,4��,
	@�6]66 0�]_[.�Y�j�	��f ��h��P2�8ɲ.��,����u	] =�P����� X���X���UQrO  s�o	�s� ���� �.�.uWY]�&�~q� xE��E��G��rJR&�P�q �+�.oX�qT�z&|�:|	|&�?D��&�����q� ��m
����W�}>Pd�&�ec�&�EX<Fh�UM�Z<L u�P<t�<H	t�<�><�du7�@8QJ/�]/+
u�
9P&�G[���'	��t���{�B`� _����
 Sx�1�zWʦ���[�_�B�� � �t"���F.�>��(un@ U�W{U��K0J�= 1���&��  Ux. t
%�_�>�'n� u��!X�.�Nl<:u(�� |�sFF��A��VR�Ђ(��r-7L+.��  �Z^�<�s<arE<zwA@($��=SW�P ��t	�.8t �PQR�e��#� �*�!ZY]� ��ECC,�&�_[�E�E��"@�v<+�<-'q�FeV�438�3�S�B�� r9 
2��������,�leڋ��+@	�	���<�YՃ� �R�
û[� [�k���H�҃�&�wU��0������t�Ft`F -�u&;Lr6A�';Tr.w(r:w �2|�	|
| ���	��ul�� bU�b$��H���X9��B�u�Ýp� ��<0r<9w,0�!��M;u	ML<u?G�	��^�@�

@G�-�2 s��ڂ��sUP��e���E �����iURV���Fa��t��G 6Bq���tW
�!u\F�\&:F	 j�RFE$�vEFKE��9@t�C&�G  t�*^"��O	O��ę:t�P�]H �^Z]�SV.�o� �<"u!C�/ r.�D�e���F�"�2���s؁� �	^[��$A�� t$?J���FC��C���s��L��{E)��6Ww>wA���_�$�L)^"��_�?z��2�)XKP��-(��\cGF��B�.�h�GC�^_XI(	P����q@!SQ���.:���AYq?RN8�r�,.�|:tA?� �����,`��O���Q�ZY��" �m�S,\8t�
3	N���$�N��<t-  )<
t%&�}r3��&�]��9q3�	C&aU:Q�Y�/�6��� ��<P[6<	t2<,t1H�u�� F:��Y&R�CM��� �\KK K8� �$� 7� ��.w;�4/u ���
� @�VS&k'P  QRWU3��޸ c�!� *��]_ZYXӨ0%i]�kBJJ
�
	 ��:r:Dw�\ ��[^D�P���X�ĴbH5�P� �t�>�	�t�n
�
'@
�	�h�L0� ��(PC�3� �$5(�S%�ʎں�% �2���Q�ZXlP� ��c�9  3ҸJ� �/�Àt	��*�:	3@��r��+)��� ���B������r����u�����ðϤ�O3�NAA���MD����X���3�Ê�k��T����u/0
�ȸ�� S������PR+�+H[ #�# P��t����U>:U�������(�:It*Du��1E���T�,��
 O��XX���� �l�%
��� �ȱ�`��}��� ���b�� &��Y6���&C �.8�=��u�;=�$�
�5"��J�WP�����VYX_�ڣ����;�&k�VQW`p�>A	�u�0� �#n2	u�� 6'�A�SV'�'$!� �-��T�
�� �PRNP��@�D��D<� �v\\�mT8Y�8G������ސ�<��hh���8�8�R\I	t0�b �  T����X%�K	 ,�a��A���L�8�82te�8 8z�8 82�_��:�:Q	,TU:z55� :�\:�U #	���&�6S	S �">�+�&� ���:��@��>���"��R� ��

�Vsu!���(u���A	�L�����8��٩� � �} '�Pp�	�S��	�S_Y|���B��K=t)p����w��>
�&e ô�!PJ��� ��#�ð	�Ds������Cze�:$�� S�8I��F��Jрt��3�A 1 ���j���`9::�*	 K*�#��0) ��P�Y�u�Le�<#�J����H
iR�?�W	�0���X �#��r'�
uJ�&�T �_+�>e��p��D(*ٹsrM�O� ��_V��B2t(�g�	X�,/* à��n E@�g�W�9��� H�=��  ���
�D� s����E����	D���� `�s
y��J��f��VQP3F(ɀ� �t$A��HJ��%����|@�� ��B �ҁ)�XY^�WV7wt	u FF���s�_;�BV�_#QV��A y� � �^(l�A��u�Y#�)VPQ�΃�!Pw$wF;�u	f�q�q��P&Z r{�bY�DX|7�>&P!t� ��,� �Pt	��&�v	XY���#h�`������XQ�Q�t`	� ��ua_(4��3�Sh�0L�Q�4G  ���������4�uN�r"�b�s_�	�Cu�NsL�ͅu ��\�hs��,-�Ih%�&8H6�u'( ^w^�� 	
;�	w	��	�	v �I?���2����w��8MY��}X(��L�n?�sP� �+�t
�ӈ8��r
���4�YN΀�r� �p�����!���?x�B��;��ڋp ��ûB	+)c	�J&�*� ���!\�83�B	:g��Bh�r���s ed�'�3��S�[ �  \�>��"��
��S�� �3����C�4��	��rlu
�1���~r�X�A7����s�G����K��Ȁt?�I���sP�����m�v�PP�9��)� I^=t���R��	;HX)�s8+"����5�4/G� ����d���,�!t�ئ���H�B�o���"���p���Yd�:m? ���,(�l���dci�*|�	 �@��
�$����P)n��" á	BRI��-/?TA��S� 6�
�t@P3Ҁ�
��X+��P����&��@�[��68T!�ȡXE��;�v�PD|Ly�[�]I70`�k%��
�|0��� �����f���a��P�M�I�u0eNu)]�P܀	�(��/
 BVu�� )�)����$ ���s"�
�*��L��m	��� G����� ,A���@��6�0��
��7(4 �C���N������]��B��Ëȋ�3���  á�
��
�
�� H�� 1
��� ����6�
�Q�O��
��1��dC/�
$���WQY�� U@ OZ��2�	 �c1��&����� ���z�4%HF(FF�s  ����
 ������=� pw#�u�^��6�u�  *�u�I�=H('w(��y(&�� !�Pٻ �����X�`����
s��HO�%%fHD���?1
��Q�b��� �	݉��� �1
 �a���&ܶ
P �� t*@vQ�@  P�SXYr�'�  J�ރ�@��@�;�3����P�ƻ us�� c ��؎ۋ� ���R�P�Z�O�����a#5h ��X�[�RTĺ�2޴�6����&�؋� �0o�}�?ء, &�� e*�����aHo�t(9����a��� ������#E�]=a�/��Q��q�f&�g�X&��T�&�jD%;���T��#�6��vF'G<!.�n'3Q�t�^Y5�؅r^4YD�6	&�l���Ɏ{��1L$ �I&;�w'�v�q��r&$"]�2�FK#l&+a�u�GL� ?���a*�Ya>u� E����R��cw	s(��n��� ���s	Z ����h��x��>t�BR�yP`&��P�R�uK.�JU.".2.�(8�G���ʟu��`/���ssgu"�=`9����a�X��r��~�C���q� ��,�	�R-/��?A� j� ���	�����N � s���>n(t
{���r�P(�:-��3�[t<�p 0 s�,�.:��@K��wu)N�-�&�)S	Q��w����������sla�/	��؝�:���U�nC�
7���7F�N$��
9 ����
Ћda�p���Q�  
�vY�B�@���3Ɋ3df>'2,!�������Sb���
�[r&X��M���WV�"5IT^P&|&�&Q)8.N��X&�{�̵�z� �r�BzId)������&PD�pQU���D<�t@�D ht8���";�Ir*B8m�ǲ(����TY �*I;�r�^Y@a�� ��
_�&X��"D.�@��� ��`�&�n��$� ����؎��V��3���6F+������_�ADx��W�@L��]��s����)�#j����=%ƒ�8fx2�<Õ����>� C��f� ����>H_u��ltu%�N���P�+�������C�+�*85 ����� ������2��ᣔ���)ҍ� �R(��,���pu	�uR��oy/ړU�	� Y�����SI�i�NU��@,�%Z��6�$:8& 8PRS�L ��r�3۱"���9�U 0������Z[+���!!+��)�� [3��6�K��A4��bQ$���̓�y2����ZP���D�l���
%A�l�`�t	1���c�(�(F
}��V�8���	!����~�p$' ��$_�F�q�}E����,$Y��~3ҍ�Xq[�s��Z��=U���uK�N05�Y��Hf��'�:3��3~��2Ѕ7v�vl0�����dG��,�V@�0뮁W(��>�Nw2<tl��*d*,tL��]zuS& 	���l��w�\��Pa(u&f_	t�9uߎ�1\�')�=���
( �C�s�����%� �;tCC������ ��>�
���"��� ����\
?��q����
���9;��Y���1�p�B3B,��Pu%�uVWQ��َ��v6��o�Y_^��^��
���&"�5���@dV��
��TyR3�Zj�e)����� @��S�
� �ɢ Ɓ��t�D;(�EuuMRr�
���U0�
�/Ҩ�:V��bU���G�p�#| �;��YQ/)��#)��)�	�A#Iޯ~ߘ���7�c1� f������\s u�9�q���l%t�X@�)t+ӱ�����u9���u7@u���i"lH0���(]�w$u\&$ �t�(��M�Y�q����uN<Ã>w��uQcw�1�������Ѩ�Q,V�>y�6q��	�ڹ�s"��u�#J��zPk����P
��L�>��D��B �@qu,���hb �2���F�����r��d�	Pz�E*`�*:�,��Z @£�����Y���q�� ?D� �#``�� r���u ��q� � � ��  ��A	�  � ���2���
  Non-System disk NTorerr Replace and pH(ress
y keP(when ady&\ ����H�
�<���ع��R V�>�@Vj{�> �y' p��T�W�C����	Fr�8����ë� f ���s���8���G��P��/�0ݑ�020UL�) �WV�ގƿ��
9�^_���ft�Go(HX���r���I=P�/��  
r`�>�U�uOw���?k9���r!�A ���G���9� �oڤP!�����4H뾺��Zm1	Q	�%� w�W��XE��X�,l���
�; 8�����Մ�1�����U�^� cÉ��a܌�A����"���F���������Jt���k ˢ�%�6�P5�r	����/���5��`T�Í>I�x������k�����I��ve%�y܎�,H��;u�P` ��%0i�-��Z�4Zo�mg�ok� GcFO�(5����2�P? r�X�(A��d�� ú�O�&�� `Z�E�G��	�-.���
����3��r�������	Q ���&��9
�؉�V�������� ��Ck���Na��	� "�H�:! �j�&�
;�v�E �SvR���g k	��	�o<S�tQ�
��1v`���t���L�n�?P�R���GC@[<Au��x��3� �*sI�[)� 
����&�?�>*u�}��I��C!q|CuD�8ZR�>(���$H�Z�ZP ����
O�Ӻ�kM��
���z��~�C1F��=�
P�esf�&d!��u��@����M.�F�(���0��V�s��(�V~i֝s�uv���]�GR���6�� sׄ1p)�Rl:9:��:�N/ :��5�Q	����u�P��
� <�>�
�J�@����C$aݪb���FC�h��؂��
8�s	<  u-�+ �ݠ�8�	|  2����؁��}�J�7�t
c�=�8����cէ���j7���àȾ��-;l�-�z�}=$ ��>�ti�yБ�7��O3Ҍ�z��s���^����&�dr1�?�t �u��u���ab�p�r�` ��&QH̌ ��S�� (�? u>�g�u�o,R�� $�r?EQw"
�0&� w6�y[�U�b=�O���T���\��L��B�
&�Ć=(��g&��8�� �|&)t�(&�(���u��������r!a �3���*����6���+��Ww���E\�Ҧ����2�R �\� ����
�.�
�%�v��:`4'����� �mt�s�E�1��,XA�;(�w;Dv��U�*�R
 6j��+�Z��J-e��>)7z3��Qz�B+����FK���!�H�2.�d���y�HxweU]N],�
�\��-]rn��+(  ?�=�r
/�����U3.ɘZ�2�(�0�*���!����"6+����X�.B�����+�iB2�a;�s��=��w�Ԡ�UX� ���؍�8QUV�2f@��!��D
�S^c;]X�� ���	R���}r��RB�rЍ��5�Y\	�� s��/s�T��⦂0�r�B)�gW�
�uU;��7�����£
�b)-�2)���8� ʉ��������K���]�vY&Yw{,��7$�:���<$�n���Z���?L� B��Fb�'���� ��=aʪLR�CQ��qD���R�%u W�H����D�y�����L����a � �O���Q�WS�YUE)�G�7�W���)2�� ���!�� r��s�;�:��` ��P�D��X�3�È�*�W��>XF}D2R��"��V�'B��K��@��_Ft�@�P�&P� ��e�����/�ft]_��;Q� �R����T��9��Ϛ�@�����w�h^��;��)f�WP)`?A��g�-d�� �=��=�tG3X�Z��w=?=�=!�=�|= leLKu�&-��`Ě����3��-���^��-�-��Ƽ�&R�����4�D(	���C U�r8�6 J��FWp  s�(���U�s�P�@>�rZ� X�r�) 'W���Q�A������Y�=A3/�x6�}le�Q1�P�~�>UQ	;S(�v��XU� 
�
Z��B$�s�Y3��!=C9;�0�Pr��$��	b�j� 2h��RQPWV�^�Y�UW����d��Ӌ>�Y6W`�

����Pp������t ��H�5I��t��ߣ��@h�^��_XYZ7*e�Ļ+�h�������0u����$q##f��
Ch�
�Eu�
  ��I����W�W,IR=L�&$`W�U@H��.Y�5,V}���'st�4�
D!�w�ڲ� ����	ö���#�4��Z���,�PM�N2;$T�w_QNP'u�F�(�L� 0����
���� �� C�a�v��!YQK�>�_< YRPQ�3�Ή����Y�FP��B�00[I��)���P`R��u�"t8P���H�)�s��"R�S�  ڌ�����������Y������5��3�$�:7*�� *�&�#� ,��&!&	;�-_��P �����@�I��ţE)�� �\
@Z���a��QWV��ϡ�ƗOצ��̠֋�z�^_k%Y�VWR'51� NG��r�+ىs����PB�G	;�@�v
͕�B���	1X�S�IR�ы�[��(�׋�% ʆZXV3�,3�w%��*��c���� 0�s�r�Ƌ����8@�	>�����*Ջ���O౑7�� �b�y�&�8��I"����&���	P �w r3�8�u��U0 ,u�ˏS�s�]7�J� � v���A�F u��t�����y�&��`+�&��&���(�&�}c�&��ROeO!|�狸+�������`�`��� �Î����t ���H��Dx�RS�r��&�u 	% �����!#%����Sm%pO���w���Uu���ja)�����r��2�'�u�}\Fw3�E	�!��C�	��,P�,�Xoh<����$�Q�8���R��s��� �/�r:�8 ��� ;�"Q�@r�@ A�( �XYrd�� ��X  ��@��@w��
��#F��� 8���
����Īa���
I�>u��	 �����PSR�o�[3	XP3��bX@?#v� #
Copyright (�C) 1987-90   Central Poi	  @Software, Inc. ��8
$<0?teS@� image % thKs�b/a.)DOS vPersio*mu ��b%2.0�:�h|% 'T<MIRROR coƢmm�c��no0�$��k@a ne*T�:k d�uU:procK�s&:ucful'u݄n)D[ x $����y3��4ed�%ingEX�t:Ttes wZt�t ���<file'E }�ckF���. C��Bn/I�"	fciP��{pfv9fofЧclosegfm*e�y3o�x8�ll����|5 Y�bod��ac.r�is��(

27�t
�ibo wi/��R#�
�4ol'��rei��� 'i!�va&a�ziir��dir��%e��  De�+�uJ�'If9m	gA�#Da}hi�d ��G�updF�Q�l �op�1��%buUit�E`loc`dU��l25 ����Ң;�a�� Ih-$=wah��ddu,�	�\�3w�Knl|u7'�DKfl;ounya�+�i�ap*�}js!�`�a���_ `�.�oX.�J��kX ��l=PPu P.�uX@��A.�P@�� ���Z�3�2@t�r�Æ���0�X��=�R#�u�)i$ W�@u%��/��   �M�� ��u�&�  $�<Nu��� �qGx�[A3�B`�S�	U.�>A�H s�SM(��T葌^�lc�h$����"r�
�
&���DT>���=Q(��oU�>qEt�IJӂ�	 ����,��.�&�X3��5��x�vX�#&�|zX�T�1Z$%))	8	#	ë W.W.�g�1
,��~X��#VWVU�� ��O�'����IU���v0~����
���0�OT��'���T '����]24Y[X��p��x:\tu.BAK  ա$FIL g!BWVSAVu�X')ܻ�0�_�=0 @�aMSESLIFVASR�IMAEP
A���� ����/��u�=1u�%��E7�6�Z����Z ��I</t ��Ar�<Zw�.�)"�"�3�U>Uu��.FQn�����"�))��V[J9nTe&e��d��fb��TT� �5��s  �S��Ss�w�2t1)u��
pXUr�����w
s]>kXP\u��87#,�O�C�!/�s�UE�lE� =C�����"FK�B'� �.�6��Z��;���r�#��KS�|t� �6�+
B�)��Z�D.���	�ō՞TrGIrB.�(�&	VP�����
�(��Ў�X�(4�EqMŌs��)������GF�Gc�p��r���-嶿S�=�)��HE���I.���Teټ�����c��*ni[^)�V��[O����*� �+��,C��QZ�>q�# ���Yt��.�It�.�����`���$G�yc[�V[C%�6W\��_ =��R������4�-��|T1?�P~[���~�����[�����"k3�)L+|�K;�8�t�7��uY+'`r��rÙ��+����R��Z� �����A<�v��B��غ�q���#�%	;v�\q�)�!�ȼ*���u
F u�t~f� t� ���2�U �2�.� [���K3���r@����xmX����""��M�@t!@��SC��'�`rBB3$ �3�	�Z ;�vO+g��O�2 2(2�*2��r�	�j��@�6 ;�)�r�]���b���L0�������C�[�R'4	 �u�6q[�  d�f[qat�SQUq`�Ql��qsX6������Q�� @���&��&­� ]�]G����= rhU�UU.��`�xI[�u2���Q$��O��	�ŏ	� }�'��Dw' ��l@(=�s#��2�'��K�3�p E�!�������~�1�hA� ؃�: 	���Z�� ����[��R�J[���LNP�4RT����<rr�Z�ZZ��Z�� A��[w���r�'K'�A '�Z�\��Z���L>)� ��Z����/-�GW4��G3���GE����U�
u��i��qr�C
4bvih��3a� 	���,�35k	,�-�Y_�@�~��p������������bH�@3�<�@�>xL)�nǺL�h���QR��r
wZY�!�*:#.V�G�/�Gq ��uL�G.: [uB�R�8R�
�G�*���G.�[�X[b�Z (މDZ��Zr�U��^�I�.#�e3�R��[Z%)�*�MoIM�$AR�.44
A�t�ؚ�c'[����O`�XU�k�p@�.��d r+3��*
��t#�����A� C�	��� u;�6�*P)%�1����
�#���t�$������A,@&���tWcAR��äVR(V��2�2�<.�O��G8@[R�� P9��ZZ�GJ������� c�[*"�[��I[.�G�v+�z Rs1�O�[+O)L�� LI�[WHY�Z��e�� ��Z�, 1��1�..��ZGz:?�%0b�*X�'��[�(s��sN
$�Hw*��X�D!�XtDs �� ʅXJ�T�K�@r�B�d<J�C�	q�Q�c�*X@�><����w+�?KC 
�D�Z���ՉD��`{�#�ZE�D� sӋ`����~w?��������Ǘ�bT��Zv��r��D6�[��  ��Z��Í�U��%qT��O-�Ou�#O	��k� U+Tf[���q<p#�õ��
$Z��R��\�J.+	w�+9k �aW���Z���Q<X,/�V��C4�C[�,�t'6��	$�A��A���"9bt\j�4����H;��{.(� * ⨧[�-�#��Q�A4���@�
3� (������8a*<��~(HE![�r~d�A��B	s�.�(��[FV�7'ɺV���@��?�t&~!��
J���=w� �Ã��(�,6)Z  �]�u�u� ,u� 8 �<�+	t>!��E�����Z
bQB z�PLJskPJsYr-�0�����O��a)���ÿ\T����H![uz|�@v�?�` ]! ��eb����� ����bc�u0R@t"Ne1>1���i���*HC�C�U
X�P���S-ͷ�#���[����[�Iу�Ji%q��@R�L[th��*
H5T[r#P.+&A.��RJ��N,UP ����T�RKtj���<RC*J:\��� ��J�������^�/tw+�� �<;��U:�f�Y�tmw����R�p�T�u`̀�*7TBwM�
76J�wA
.
;9P<9A�yh�; z��������b��PC	����47r��I�u�UE�g
s)�S>�6�!���S`X�ė�>��`c �i���@:Rfd8�5��q���?U�	f;�r8H���A���D�i��m�%�Wt�D�Z�.r}�A��
�s �Y�Z�Vo{�\rr�=�'&wB�����
�Z�He5W�<<��YU4U�EK
]�{tv�� X2X��X|9Xu>WU.��6l�Z�A� ����1ʜ���R@���Zv�ʌ�)@ T,A^EB?��t��
���%r,�.� �K .�9 "$4��5j7+]�Ý���jPQS�آ�<�{[����^ ����� ;t��r%�&r
���� e.����1�3��J�+=�J��� ��?�s3� � ��n��p�*	7�;�&
v0�63���t��CrQʸT ���������O�6	���/�/� �PR���ZXtEof#`t�9Qjj-�(�:+��l%,Rl�=��0 ll!뒥;-ggU$*}*xR�x�j<j���Lm)m5m�4�m+m.��@m5m�,RC�:m��` m1m3�$�Jw. n-nJ	++�k��3��h��i;iGi
�i=i����@!r��6?l>A+>#6����xP ��-
�}�F��LCu ����6H�>J�Rh>�)��PUe�R��(<yg&t^�(/$�5�^��u:�b^� Ju�  !N����(;N�{�:�^xvx�'x%� ���.ti�  x x*ۦx)xx1mzx3xu�x1x� xn��x� 9x7� �>��gu7�	A�o��r���T^>K>I F ���7� ���<�!���r�ϋ��3n3ɴ�j�� ��= u���ڣ����|*銻�Äbl:NuD���X�o� ы�>�^��  r�>�F>;Fu
�	v�u�4t�>�FH�3�r�>�^ 7V���$R�Zv  +��WV���� � ����^_;pv	���T`�J|�s�E����t��V
�=���o�
���� ����� �> t9��t	�fh;�h)B\	>T�5��v�@�@����N@�@@�]@@%�@@@%t�@'@ �)@�@)@f�n@+@+@�J)@@-J�@/@7@96�@�@�?r�&r�;La% 6?��6A6I6Kk6�&Fǋ�i`4��� `L�������Pz�!�X�PRU�� ?�]Z(@��X������u���6��_ ����E�����K  �Q3��t�6�+�!���. �+�m	�Y�ΌQY���l$���
���
R1oP0����XZ�� ��� X�i��&�3����v��
 ��u� ��
P�t���
uD ��ږV� ����r-Y����;���K% �a 
^���@ 8X �u���s�^+�Ot:�t  ���V�ذ\&:E�t��&��&uu�
��u�^��0VP��H��N\rU7Q�Yu�C�� �E J	~Sp<t	.O@���Ɇ!t �]BAo�bO�.�CI�O���]  iW� ����� ���-O� �	*"G�<�ǧ�Bu�z���QH:_Í6U�L9�6P@	;�3�&�E, ���VQ�Z^tO2(�� S&�=m�|�u����
[P���lȉO�	&	E)�	 �	 $��>(�� ~��&�P����&. ��7�����o��� ��+@��X��WYg���o ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  �Y                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       ����  ����  ����  ����                                               bc  � 2@          22                                      � em  0 ��������������������������������������������������������������������������������                                                                                � ��� w                            I         � �   �����    5      �8�=   �,�+�+� ($�" #"#M#�!�!Y#J$�$�%�$�$�$�$�" $�"�%�% &�"�++&O&�&�&�&�&�&B(�)�) **�*�* +!+W+x+�+:,O,�+�,,..�./00                @ ` � � � �  @�� @�� @��� �   P  @                               �?������  ?  ���0���   @ ` p x | ~ � | l F     �?������  ?  ���0���   @ ` p x | ~ � | l F     ���                    ���   @ ` p x | ~ � | l F     ���                    ���            �                                                                                                                                                                                                                                         !   �	
 !"#$&0@t~@ABCDE`abcdefghij`anopqrxyz{"#$'(               �  �  �    
    X                                                                                           		%')+	!%).	#'+05< $(,0 $(,048<@ $(,048<@DHLPTX\`                                                                                                                                                                                                                                                                                                                                                                                                          	#(,159>BFKOSW[`dhlptx|�������������������������������������������������������������*** This is Copyright 1983-1992 Microsoft *** �   l �#, \)� �/G 05 x           �               �   �                                                                                                                                                                                                                              �I�I>J[J�J�JK�K1L1L#L��� ��� ���	 ��� ��� �	 �
 �                                                                                                                                R  �G *** This is copyright 1984 Microsoft ***  �?������  ?  ���0���   @ ` p x | ~ � | l F                       ��  �?�F������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                           ��������������������������������                                    �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������s�������u�� ���7���3�8mu�8Mt8Cu�L�L:Mrƈ&L�C�>; t��6�tM������8Ù�>3�8�+�l*��S*�8��t�>> t�>:t�>7 t�����<+N���F������:���>5�:�-�-*��*�:��t�>> t�>7 t�����>+P�Ȼ�?t�?t	� R�1�Z�>; tH�>9 tA�>8 u4�<+N�ŀt���ǀt���9@w��؎��9�8���r�%	�>�<�C
�t52�8&nu-�nP�[$�t#��uXP#Dt�D�u�DV���\^�L��9XP"t�>, t�!�u�?�9X�t��E�m
u
�����m�nˋÌڎ��G >�2��R���.O����S��׿ ���S�؋�Z���.Q����U��׿ ���U����PQ���y���y��;�s���>�2���O�s���I��YX��3�8�t�9Jt�S���.T����L����>X�L�؋��.V����R����>X�R+�X�.V����P����>X�P��.T����N����>X�N��3���&�$t��s�����Ȣ[�2��P�<8>vt����>�6��>��D�>�^ �X���D������U��W�v��v��v��v�<+t1<.t-<	t9<t-<t1<t%<t)<t%<t<u!��T�|�t��������t����ߎ�PPSQRWVU�^���]^_ZY[X�~��~��~��~�X<,t<-t<t<t<)u�~���~��~�5��v�_]ˀ>. tv�<�>v t���лo�?r
�?t�?u����=�v���>2�С>���>(� v���>4���&P����t����̈f�^�n�V
ˀ�t���u<0u�F�ˀ>= t��r

�u�8&ru�UP��2�E�X]�F��F��I�F�ˌ�3��ؠI$��P�@<t�A�:t"���<�;�?�>�2�8Bt��;�>X8&>t�q3�"�o8&=t
P�F��SXr
�~�t:t��b2��)&�ގƾX����&ˀ�Su	P�/ �3X�)<t*<u!��u���uI�N���N�ɉN�A�N��F���F���F�ˉz�|�ێûx�^�F ˀ>; t2�>< t+�<u%��؎�������0 �8 ������<6s<.u��2�S����؋��[���<Mu�ߎǿ��<mu�ߎǿ��Hu8�D�+�-����+<+><>�D ���C�q �P����Hu�D8Eu%�� Hu�>D u�D�8Eu�m�D�m�R���������&3����������&5��8  �:  �<�>Z��A �t�������A �t��� ��t����A�t�
����F �2���4 w�o�>r u<�>>u�� �-��D��D$�>> t�61� �>>u��P�Xt�0�o�>w u�)�2��7�>; t��.���>> t
�����B����3 �5 �&H�/�(H�13��m�n�S�U�,� �ߎǿ��P�@�B�sH�E8wu�w������0 2��l#�>; t�F,�X.��	�X�����L#���&�(�����s�ڊ�3��ؠV��<@t
<t��ð#ð&�;�|�ʀ>v t��������/�>; t�z*�;�|�ʉ�1�>; t�E*��+�-���y"�؋��h"��+�-�>> t�>:u�>v t$$�� �>7 t��>8�.8�>> u	�>v t$��<�À>> t�>:t�>7 t	��>:�.:�>�>; t�.3��8�:�8Eu�m��m���ی��؎Ë�����2&8;t�B�[�#&8>t	��� ����3��(8;t��*��,3�룻E��?�u����P2�F8&v�<t$��F�>��F
þ��t�3�8v���F�Dt$��F�D�F
�P��Fþ��tվ
�Ѐ>; t�T-���E���Ǌ��壌�>��.�����B��Ø�>> t�>:u�8��t�����@2��8!�Î��޿��  ��� ��� ���ؾ��� 󥾘�>: t'� ���>:u�$��� ���2��� �)�>8 t���Z��� ��F���?�2��8Et�>E�u�m��m�E�2�8;ub�E�78>t�u�X5�;��-�+��t8lt���� w�2�4���u
�t@s�t��E�"�"Ԋ�ʴ�D��D�3�����F3�����F
��.���. ��uA�uB�3�5À>v t�>> u�����������7�9�6;�>=� �8.Eu���>�<�8:t8.>u�8.7u���2J��4I�28.>t8.�u�+B+@8.vt����BB������JӋ�ZI�Ds�>D t�>; t�C+�m�o�m���<�>+N+P��t��E�z��?�F
�A�F �2�F�A��?������? �u&�> Gu
�,�!$��!á3�F����������
8;t�B�[��
8>t	��� ��
�Ë���
u��F
��F��F�3��F�F
�FH�Fød ;�r��;�r��;�r�Ћ�
��¢J�Q
�M�âY�C
�O�ƢZ�5
�Q3��S�UÀ��G�>u��	3��Y�F�Z�F�J�F
Ëãd�&b`�^ád�F���
�>u� ��D��D�/5�w�>B u8�D�!�D��;�u,;�u&�����َ��ظ/%&�D�!&�D������  �5�D�!�D��;�uA;�u;�����>� u�>>u�����َ��ظ%&�D�!&�D������  �5�D�!�D��;�u;�uf�D�����ظ%�!�����D��  �)�5�D�!�D��;�u/;�u)�)�%�D���!�D��  �>� u�>� t�F�����F ���F�>t�/���	�&*"���"&+
����z	���>� uI�>B uB�/5�D�!�D��;�u;�t'�����؎������ظ/%&�D�!�����D�>� u\�5�D�!�D��;�u;�tA����>>u�>� u������I�E�؎������۸%&�D�!�����D�>� uG�)�5�D�!�D��;�u;�t*�����؎������ش%&�)&�D�!�����D�>u�ێûi�D�� ·��D�>� uB�5�D�!�D��;�u;�t'�����؎������ظ%&�D�!�����D�/ �3�F�t�w ���3��F �2���4 w3���7H�F�>; t��%����w�WáW�Fá���F����F�VW�������5��&3&�����_^�VW������&3���_^��8 �>9 t�>; u�9�8���  ���� �x� 󥾘�>: t'��� �>:u����� �{������� �����>8 t��àG2�8&7t�>:u �F�m�F�D���F�F���F
�2�w�F�&H�F�(H�F
�3�����F3�����F
�2�F�4�Fÿ6�%���B �5:tC��É�F �r< u2��o����r�o ÿp�u�5�2����N3��F
�F á@�F�B�F2��F
�E�F��F���ǀ�s��2��࿀��%�l�F  ÈM�F  Ë��0r���u�����D�L�D ���F��Ã��u��F Ã�w>K���ڌ��؎¿<
�� �ڈ������@
��
� ������<
����N��F���3��F��@�F�^ �F<
�3ɿ�����t/K�����w&��������@
��
� ����<
���Ý3�2�@�FH�N��������@�F�^ À>� u'�����  �@���
�t	���	� �����F  ��F��ø���F����=u�фs�F  �À=u���=u��>D t�H�P�IP�-��2����JJ����>&tG�)�5�D�!�D��;�u;�t*�����؎��)�����ٴ%&�D�!�����D�-������pJJ2���hJ�`��a�����XB���Q����3Ɏ��l&��&:t��$�&�*�:�s������'���R�Q�&�*�:�s�YZ���������I��t�<����u���F  X�X��á�F��F�/�F�1�F
��2�<�>� u�0"�t"�t��u�.E�D�>� t�C�J��H �D�F�>� t*2Ҁ>C t���>B t���V
�J��F�A$<2���A$02�F����FÿJ��h;�}=��������y���Z ��*̋ي���܊���u
�t����ۨu������ۉT�Vø���F�  �F� ��F
3��F�3��F;�u
�FT�FË�����������
�Iu�� �W�It��Y�It�Z�It�J�It�����ItؠG�ItѠl�ItʠM�It�2��It�2�8@u���It���t}�J���tt�&E�E2�C��8'u��It`�&D�E2�C��8'u��ItL2�8Ct���It>��Dr8Q�<
�D�Y��Dt(�9�It!�:�It�;�It�@�It�>�It�C�I)NÌ^ �F
�Ã��u"�9�&:�F�;�&@�F�>��F
�F  À�w;��w6��dw1�� t,��dw'�� t"�9�>:�;�.@��>�<���F  Ü��-����2�8Nt�@�G
B�?u�>OtJ�G��������u�2PS3�
�t<dr�d�@@���2����؋[Xt�2 ���s���Q3����"�t"� ����D"�u��:���uY��t��Y���YûB�M�-����3Ɏ�&�l�.I�u&�l*�:�s��������:�u�>��M��� :�t��u����M�Ì؎������<
�� �����ؿ����@
��
� �&�2���<
���>��À>t�/����# �*��
��À>t�/���� "*��� � À��u<v<4w<3s<1s<$w<!r���À>; t�^<`rÓ��~ �b �2�R�j�I���>> t����t�x�83����d�v�\���>>uz��#u>� ��^�&a3��0�<�=@�:�8���.�,�&��(��4�z	c���&u:� ��^�&a3��0��&�J�.�&��(��:�8�4�U��r�M��u��آo� ��^�&a�؎�3���&8&>tS��J�6c�ǎ߉60�.�0�?�>> t�[�2�&��=P v��������(� �,  �z�=��4�:�8�&<�&=��sP�>> t�,  ��s>��s5��s�>>t 8 2�b� �>> t�4�: �(� ���&.�&:�&8�>> t�&���b ��t8�>> uQ��~t��
t���@t��tu=��~�&(�&4�0��b  ���$t�>C t�o�D��D<t����	up�&.�&&�0`��_�a�2����zG�b8&>t�t�&���&,�&.�v��8 ����R��j���@�v�,�.��>> t��@s
��w���r����_�a3��0�<�=8>u�,P ��t|�t ���u�i��\8>u(�����x:F�zkF���>�R�>�j�>��t4�(r� �v8&>u$�8 �,�.��E�RP�j��b �U�>> u�(��4�b  �>)qt9�t ��\�>> u(�����x:F�zkF����R��j`��r�>> u��em�Rpm�j�m�(^�4��tQ�>> u�b S�� � �D��D��[uU�&��>> u������t�x�8�z�=�� � �b  �>> u�(�����R��j`��4�� ��0u:�8 �&��(^�0��2	�43��b�0�<�=�Z�.�,��2�8��r�8 �>0�uq�>\ uj�>>tc����"t��u�_��a�d ��_��!t��u:�a�b �8 �&��(\�0��.Z �2	�4�<�=�(�*�>>u/�>:t(�02�U�D��D]��@����*��2�������(�&H�>v t$��/�(H�13��68t��2�78't��4�8&>t��D��D��À>C u1�>>t*��r%��v"��(w��'s
��$w��"r� ��^�&a��ø ��^�&a��
3��0��&�J�.��8�:�4�& ��#u�(��À�$u�(��À�"u�(�����t�( ���(���U��&�>> u� ������H 3�&�6��&8>t�2�1 &8>t��&�.|&����K�� �&��AA��;�r�&�Z]�&�.���&��&�>/ u&�&x�խ��Ju�&�>> t�ë��ê���V&��H&�&��؋Ȭ"@�u��&�/^��4��ϋ0���B���J��B�����؎���>D u���>; t��>�<��G�E�>:u��>> t� ��8.7t�>7 u��v�I�>> t�U����4�F �2�F�>8 u�?��>8u� �/�F   �F���4)G�2)E��4�F �2�F�2E�� �F   �F���2E�� �4�F �2�F�4G�� �2��)E�� �F   �F���4G� �4�F �2�F�2E� �F   �F���QFF�4)G�2)E� �2E�u �2E�k �4G�a �2��)E�U �4G�K �2E�A �2E�7 �2)E�4)G��]��G�E��2J��4I��	s��E��D �G�E��2J��4I�	r\�>>u
�xQ�>r t�>7 t;*s=;&s7�	�>? t�0���u���t�&����(U��#F3F]�D�hFF�+@�>> u	�>v t���D+B�F�>> t�rf�>� t��I��$��S�;��BB������JӋ�ZI��r-2��
	�k��>ot���C������E�N�G�P��E2��(8>t�Z8t��>:u�� 87u׾I�>> t�FF�>8tNN�o �>8 tg�4)P�2)N�W �2N�M �2N�C �4P�9 �2��)N�- �4P�# �2N� �2N� �2)N�4)PáP�N��2J��4I�| uFF�J��FF2�8st8?t��0���u���t������G8?t��0���u���t�����؎��2���>���>� t=�R�j�I���>> t���� �R�j�Z���>> t�b��D�6F��������.���>> t	���2�g	�&z�؎��խ#3�CCJu��"2�CGG��Ë.���D"ÿ6"�*�t>|[�����>> t��� �Ǿ��>> t�2<s�؋����G������Ȉ��u��V�َ��ȋ���2�2���
ÊܪJu�^��؊����>> t��� �Ǿ��>> t�2���N<s�����O����������u���V�َ��ȋ���2�2���
ÊܪJu�^�À>� t=�R�j�I���>> t���� �R�j�Z���>> t�b��>R�D�6F�H�6J�(��/ �ݎt�>> u�>ou�t�L�����t�]������+T�>ot������+6V�΋����@@�>ou���������6j��� �>ou������À>� t3���R�I�>> t�� ���R�Z�>> t�b� ��>R�H�6J�>> t�΋��DQS�VP�;��3ɋ.��S�>� t5�y�j��>> t�j�� �j�j��>> t�j� �4�6j�>\� �.X�6V�6T��>> u�>ou������,+��щf�.h3�Y�>> u�>ot�������}�����
f+.~
���+�Y�Y�}K�ًـ>> u�>\ u	�>o~u�&6f�������,6f��;>0r+>0����6f�����
h+(~)h~g�6h�ێ^2�>o#t8.>u!8.\t�t�����sP� ���X��u��+�t�ʐ���������ۀ>> u
;>0r+>0��uَ���;3��(8t��t38>t�@������>o#u�T�6V��6\�>> t�� � �>o#u�T�6V�b�6\�>> t�� �G� �>� t=�R�j�I���>> t���� �R�j�Z���>> t�b��>R�H�6J�����ݎt�>> u�>ou�t�7�����t�H�������� �>o~t��>� t/��j��>> t�j�� ��j��>> t�j�>j�X�0�ӡ�@@�>> u�>ou������+���,�t�݀>o#tO�>> t!�ы����6\�˃�����������u��@�>ou�6\�d����,�6\� �;�r+�����6\�m �r���vP� ���X���ø�+��X�>j�V�y�~:>�GGBu�3ۋT��y����+ڌݎt�6\���� �������y��P����ä��݃>|v�����ÿF3�>( tA�D�H;�}��>ou+�= ����+�= }�T��J+�}�؋�6Z��;�~�D$��T��V3�����V��X�T�6V� �6\À>> t��..�I�ޖ�>ot�������>o~u�x�"<2������ˊ=���..�>o#u�^ ��t�_�����64�&.�����62���3���9du&>N�^Ë6�>/�(�6�>1��6�>/������6�>1����;�|��;�~��À> t;9|;=;7|;;���À>>u�
�t� 8\t�8>u�]��=w��؎�2�H�����������^�� � �D��]	�Ļ��ċ߹	 � ��Ļ����>7 u#���ٺ ��ڸ�������B���J�Ĉ�ٻ|� �� ��D�3�8\t�8>u�]��=s��87uJ��� ��ں������3�B���J�ĸ��%�����B���J�Ĳĸ�����	�B���J�Ċ����2������������^�}	��� �D���߹ � ��߃��� ��DËխ��3ëJu�2�����Q�݋����Q�݋��������YÎt����&�����>/ u5��BU��&�%����&�%�G�CCMu�]��&�%��CGG�۰��J��&��ð�BU��&��&���&�����&��&���&��G�CCMu�]��&��&���&���CGG�뫎t��S�?��� [CFJu��>> tCF�����&���r2���s4���u�ô� ��D��Dô� ���� ���� � ��� ��D��D�3���&��&%0&��t<0u����t
��<0t���/À>@ t�SQR����,ꢒ�t�����	�t�� ��3ۜ������B��J����t���C��ٱ	�Ί������B��J����t���C��ٱ�u���<r ��t�����B숇��t����C�ԋٱ�u�����������B��J����t���C��ZY[�P��$<	t<t�X��6�&�4��`t.��@��t;��@��t3��@��t*��@��t"��@��t��@��w	��r���2�������QWS���>@ t*R�M���G(ڴ��
�t
�M���G(�V� ��^Z�_V�M��G(3����c������������< ���G�< +�������	����N�	���N��k3���
@��^3����M� �A������[_Y�����r���w,�VP��% ������7X^�
�w�8&@uV����^�F���F���I�F��P��X�3������O�� s��^Ê�^ËË���� ��MƄT��Os!2�� ���uP�u����X����������È���3��s�W����O3������s��_�W����M���A��y���ێÎ�3����Q��s���Y+��%���uP�u��Y�X����R�P���X��G@�ݝ_�3�� �W��&�5��O&�E�������_�WR����&�5ƄT��M��O&�E��&�e�$���uP�u����X������P���X������Z_�WRQS�؎��M3�8otU�o�O��w����s���+��Ŋ$���u<t)���u<t ���u�P�u����X�����P���X���F@�ȃ���m|�8.tI�.�W��	��S� �����G� ����?�u��7�>@ u�̠
���$�ʠ��[YZ_�WQ����2튍S8.@t��u��HTtI��M�I��y���ێÎ���s������Y_Ì؎���^�F �XX^�F�ˋ��������à�����>:��������>:��à�����>8��������>8���P� �8�:����������ڨu��������0�B�؊����u ���� �8�:���İ�B�u����������	�B�J��$@�ǀt��u�ࢅ��B�J����@t��&���t���H����@�	8>�u��������&H�/��B�J2�t���@t����B죐���.:����~2����1@�(3��v���������?����B�J
�t��B�t���XË�����R����Z����ú��7�B���������7 �8��9 �:?���0�@�&��@���3 �@�@�@�Ë���3�9Ft�9Fu�F�?�F#�t�= w݋F#�t�= wѺ���B��PJ2���B��PJ2���B��PJ���B��PJ����B��PJ�����ĸ�B��PJ���B��PJ��ָ�B�J��P���B�J��P� ����~�>�2��������Բְ���������&�&��θ ��v�ĸ�^��t(�N�~����������O����G����O�G������u��-�N�~������������O����G&�=���Ǫ��G������uӋ^�ְ0���@���^K@���X�X��X�X��X�X�X�X�X�Ë��3�����u��t���^�N���P�77�B�J��P����3���@����#�}+�3�@���@���1���X�X�þX�B�&��ȌߎǿD��ī����6��6B��P�DP����á�
 ����
;�wL�� ����;�w;�>�<+B+@�>v t����BB������JӋ�ZI�z�r�Z��m���R�� ��+B��+@URP����]�Ë6��>��7�6��>��>�v+6B>B������.+�>8������.-�>:����E�@�B������ �k����_�������7�B�$���������������8Ù�>3�8��o����.8����~2����h�"��>8u$�<�:���>5�:��>����.:����~2����6�"��>�<��+N+P�5�8t6��>:t87t�8�t!R�����a�P����Z�B��U�$��O�JX��Z��������BB������JӋ�ZI��� 9:t�F�.��>:�F�D�.��>8�D�98u�>v t�>D�ÜP�o�D��D$<@r��<Ew������&�X�&�$P�o�������B���X��ߋ0���P�	���B����JX�>:u�>� tN������>ow	�>ov�~����d�B���J�İ��W���S�B��N�$��>oer�>oft �>ojr`���>:u�>� t�ËL�������ꡅ�؊�A���ã,=P v	������&�(�0�?�b�4���:��2�8 �������B��
Ȁ�2���Ë���D��>d�����Dú��(�P�D�F���x��#�y���+�#�y���+ۀ� w< r� �>� t:�u	:�u������U��������0�B��+�PJ����#�B���PJ�����B���PJ����	�B���PJ�����B����P�����J������B����P2�����J������B����P2�����J�ΰ����B���P*����İ����B�JP�����B�%` ������������
��J���B�$�
��J���}�B�P��J�ǆØ��  �ˀ��ۀ� ������>^�ǿ����+���!������X������5�B���J��X�������"�B���J�Ĳ�X�������B���J�Ĳ�X�����ܜ�����B���J��X�����ܜ�����B���J��X����ܜ�����B���J��������BX���J�����BX���J�����BX���J�������BX���]��>� t���x�� �D#�y+ɋF����t��#�y+ۺ����0�B�@t��������B�@t��J�����尜�������B���J��@���ܜ���
�B���J��@����ۜ�����B���J��@����ۜ�����B���J�İ��������B���������J�X��PQ��  �ȋŰ������B���J��H�ۜ����B���J��H�ۜ����B���J��H�~ۜ���x�B���J����YX#�tbPP���"�t �ŋŬ�����Ŝ���K�B���J��H�ņ���"�t"���$N���Ŝ���)�B���J��H���Ȋ���u�*����"�tFXHu�XÜ��������B����PJ������B����P2�����J������B����P2�����J�����B����P���J�����P����B���P*����J����B���P*����J����B���P*���y�J���r�B��m�P$���f�J���_�B��Z�P���İ���N�B�JP����D�B�%` ������������
��J��*�B�$�
��J����B�P��� ����� ��X��������B���J��X���������B���J�Ĳΰ����BX����J�����BX����J�����BX���J����BX���J����BX���JX��X���ٜ����B���J��X����ٜ���y�B���J��X����iٜ���c�B���J��X���Sٜ���M�B���J�ĝòĀ>ow�>ov������ �2���� ������ �2���U��ދ�������B���J�Ĺ  ��������K��s�]ú������آ�����B��J��؜�����B���J�İ���B�� J�؜����B���J�İ�����B��آ$�Ü�����&����p�B���J�İ�&�_؜���Y�B���J�İ�&�H؜���B�B���J�Ġ�þX
�u:
�t63�������ߎ؋����-�� ��ؿ��&�E �ЪG�������u����؎��?�3������������      9L ��  ����  �     �k�k�kl�k�k�kll�kFlRl[lkl}l�l�k�l�l�k�k�l�k�k�l�l �(C�I~�_2E6(5�5p3K6.5�5�2}4���� ��� �,�2���!A(AZC`C  ) < j ��#%�ld�!�35�!���t��3ɺHT�¸ �3�ǁ�HTu;ל�3�tw�ǁ�HTuo;�uk� Z�6Z�4Z�# ����3���t�W�� �� 3�
�t�9� re
��ug� �>3Z t��>(Z u� �  �3�$Z�u�$Z� ���
�=+�� �� 
�t[��� r�u'�m�u�$ �$Z�|�$Z�t�$Z
�l�M�(�$Z�_  u\z\\�\R]�]V^[^`^e^#3C"2B�/�+P� o3����PHXu�C� ��؀>���u6�&iZ3ۺ �%Zt���[SR��Z[s2�>�[ u$����� v��%Z �u�%Z����[ �$Z��[���&%Z�9%Zt/�>%Zt(���@��s�QV��[���%Z&�� PW�FJ��^Y��>��:��6��2�<�t�<�t���ع �<�u��:�u���OJJ�-�! ����r
�t"��uY�>iZ tR��/��I��[
 �$Z��8iZt)�1��� �/���r�
�t����	u�1 ����[ �$Z�ø<+-��������v��h���)�Ո.*���-�ú?����԰���JJ��԰BB���JJ���:�t3���B��'2��l��2�
�����
�u"P� ��؀>���Xu��#��[ �$Z�I���u���uA��uA���)� �*����-<�>���ହ%�ô��
�uU&�G�q<�t�t<�t<�w?�)�0�!<r3��t-��>�㯹���-�)�,)~�)rZ�Mf)Y))����þZ��Z��Z��Z�� ��H��Is"��H�.H��I�.I� ��H��IsÁ�Z����Ƣ����������@�P�-����5Ӱ��/�B��R�/��#Ӱ
J���Z��
 ����R�1���Z"�2�"�t/�����R�1�Z"�"�t�ӊ݊����s��C����u�Ȋ���2����R�1���ZXR�/�Z��V����-��)��*�-�����P�����JJ���P2����J���P�`�{�����r��JJ�l��P2��e���aҀ��[��J�V��P�K �-s.X���X���?��BB���7���X�/��BX�)��BBX�"��^��B���
���),�^ð����3��ػl��:t�.�&H�*�:�s�����J������ьʎº ���v�$Z����+�QWV��+Ǿ�Z� ��=t
�=u��Z��<FF��^_Y�>D��s���"Z�D�ȣ�������������������������,����D���)�5�!����� ��ؿ�?�����4�xV�9��t � ��ظOL9J�t9P�t9�t9L�u6�&?�Ȏ��y�>>u�ߎǿ�D�>�2�	c� ���"ZE�� �e��0� � 3���u� � ����Au� �>�"Z�?�Du��G� ����ͫu�=��3��
߈�u^�"Z�?�Gu�9L��7��3�8>t�3 �j��R�8;t�3[�>Bv	�@�>�;�؊&I�c�ˎ������ 03ɋ���t�>�Ȏ��@ �&W����	� � 8=u���u�������Tϸ5�!�>� u�>>u�������I��������/5�!�����35�!�����5�!�����>; t�>��6��6B��P�XP�`��� �>0Z t�" �>N t��ȣ���R�hZ�=�, �I�!� K�>�!�u��&3��3�u�&� �$Z��&���"Z�'��L�$Z�!�t�խ&#3�CCJu��&"2�CGG����ۀ>~ tP�ǀ� |'��@|��`}��  ���  X��ۀ>~ tP��H��X��݀>~ t"P���@�� |��@|��`}܁�  �ց�  X��݀>~ t�P��H�ԋ�+D��xz�����������������������>� t����¾��9 FF���7�FF���jZ��FF���6D�"Z+���s��Ì؎�2���8>u$�B��` 8;u�Z�>>u�78�u��
R�@�Z"ZD�ϸ 3��<u?�B��t��u����t��t
��t��u�@�A�>@ u� �>; u� ��p t%���
�ue&�Gt^��� ��������K uH����2��B���$�<u4�;�<�"ZoQ�>� t��B����` ���B����` Ë��������������������ø o���7Vu0�>�?�"ZZ�>� t�������X������ø �3����KOu�>ø ���&�>��PuA�����t8��t3�ߎǿ�D�(c�= ���Z��D��Z�譋��ª��+ǫCC���"ZfEú�������2�
�x����>áW���拴��RV��	�!^Z��	�!ù` � �3��~t�� � �3��� t�� � �3��� u� �$Z��3ɸ �3���3�  �u1��3� = u-� Z=\ u%�ӌ��ظ3%�!�ʎڎZ�I�!� �f��$Z�^��$Z�V��&.�D.�FU��L.����D].�D.�F� .�D.�F<.t
�u�PSQRWVU��L�U��]D�.�>� t.�D.�F.�.�.�D.�F�.�D.�FPSQRWVU����^��U��]��d��.�D.�F�.�.�=Su��vW��r�P��uK<t<uC.�D.�FPSQRWVU����^���F� ���~� te�~�u'�����.�D.�F�.�>� u.�>� tS.�.�.�>� u.�>� tU�����.�D.��.�D]���^��v�������]^_ZY[X.�D.�F�.�D.�F
�tO��tJ.�>= t���t=��u<0u4.�>� t���r���v"
�v.�D.�F.�.�.�D.�F.�.�PSQRWVU���
�^�U��F�  ���~� u���f��>� tR��� ���~� u�^��,��� ��.��U����� �^�^�~�u�v������~�u��v�������� ��.��U���� �^�^����U����F��
U����F� .�D.�FPSQRWVU����^���F� U��]�~� t%U��F ��.�D.��.�D]�^��v�������]^_ZY[X.�D.�F�~� u��]σ�]ˋF�^�N�V
�~�v�F s�^�nÉF�^�N�V
�~�v�^�F ø
�/�t� �/�u	��F�/�u3�t� ÌߎǾ�f�\ �׹�����3%�!�����%�!����/%�!�����)�%�!�� ���%�!�2�</tG$�<Ou��t�$�<Fu��t�$�<Fu�3Z�(Z��u�2�83Zt8'Zu�Ё>%Z��t@8(Z����*��ՠ)Z"*Z"+Z<�t2�����J�Y�Z脻�,Z
�x2�����>1Z t����3�84Zt�81Zt�03��3�J�0�3�>2Z t3ɸ0 �3�D�C�0 �3�>l t	�.Z�.�3�/Z
�x�.�3�)Z"*Z"+Z<�t)� �3��8)Zt�)Z8*Zt�*Z8+Zt�+Z��3�,Z
�x2�� �3�W�" �3�Ύư@�&Wۋ�. � �3�-Z
�t2��- �3�Q��3Z%� �؀�A��w����5ZY����0Z���'Z���u��%Z����t�= w�
�t��%Z  �&%Z��u��%Z ����+Z�J���)Z�Y��� t�= w�
�t��%Z �&%Z��u��.%Z�%Z ���DrX�2Z�u��� �W�l��l� u�Ǣ.Z�\��z 
�t���/Z�M�J��h �J�1Z�=��[ �t= w�-ZH�����$��+��? u�$�,Z���e �*Z�Z�U��Y �*Z�Z���� u��@����� u��%Z ����QR3ɋ���Ǹ
 ����s���u��؀�0r��	v�N��
�ZYù�������u�2 =d v�d �Q2���O ��<Ft+��<Nt+��<Dt��<St*����<Et��<Pt��<It2���N�Ǌ�Y���� <Lt����
 <Fu�������<ar, �QR3Ҋ�6C��Ŋ�$�<Pu�C�taH= s[�S2��؁�F
7[��<Su�$�tBH= s<�S2��؁�F
[�<Cu��u#�.C몀� t���/uN�����t��
t2�����̈́�u�
�t�6E
�t�D���ZY�MOUSE.INI MOUSE=EnglishFrenchDutchGermanSwedishFinnishSpanish
PortugueseItalian #o�p9n�p�p�p�p'q;qWq�r9n�r�rs*s[sos�s u9nu-uGu^u�u�u�u4w9nOwaw{w�w�w�w�why9n�y�y�y�y�yz'z�{9n�{�{�{�{+|?|[|�}9n�}�}~.~_~s~�~�9n�1�K�b�����À8�9nS�e����ǂۂ	MouseTypeLanguageHorizontalSensitivityVerticalSensitivityDoubleThresholdActiveAccelerationProfileInterruptRateCursorDisplayDelayMemoryHardwareCursorSupportForceDefaultCursorRotationAnglePrimaryButtonSecondaryButton	ClickLock[AccelerationProfile1][AccelerationProfile2][AccelerationProfile3][AccelerationProfile4][DOSPointer][WindowsPointer]PhoenixBIOS BusSerialInportPS2MSX LowMemHiMemEMM FalseTrueOffOnNoYes LabelMovementFactor PointerSizePointerColorGrowth	ThresholdDelay SmallMediumLarge NormalReverseTransparent 	MouseTypeLanguageHorizontalSensitivityVerticalSensitivityDoubleThresholdActiveAccelerationProfileInterruptRateCursorDisplayDelayMemoryHardwareCursorSupportForceDefaultCursorRotationAnglePrimaryButtonSecondaryButton	ClickLock[AccelerationProfile1][AccelerationProfile2][AccelerationProfile3][AccelerationProfile4][DOSPointer][WindowsPointer]PhoenixBIOS BusSerialInportPS2MSX LowMemHiMemEMM FalseTrueOffOnNoYes LabelMovementFactor PointerSizePointerColorGrowth	ThresholdDelay SmallMediumLarge NormalReverseTransparent 	MouseTypeLanguageHorizontalSensitivityVerticalSensitivityDoubleThresholdActiveAccelerationProfileInterruptRateCursorDisplayDelayMemoryHardwareCursorSupportForceDefaultCursorRotationAnglePrimaryButtonSecondaryButton	ClickLock[AccelerationProfile1][AccelerationProfile2][AccelerationProfile3][AccelerationProfile4][DOSPointer][WindowsPointer]PhoenixBIOS BusSerialInportPS2MSX LowMemHiMemEMM FalseTrueOffOnNoYes LabelMovementFactor PointerSizePointerColorGrowth	ThresholdDelay SmallMediumLarge NormalReverseTransparent 	MouseTypeLanguageHorizontalSensitivityVerticalSensitivityDoubleThresholdActiveAccelerationProfileInterruptRateCursorDisplayDelayMemoryHardwareCursorSupportForceDefaultCursorRotationAnglePrimaryButtonSecondaryButton	ClickLock[AccelerationProfile1][AccelerationProfile2][AccelerationProfile3][AccelerationProfile4][DOSPointer][WindowsPointer]PhoenixBIOS BusSerialInportPS2MSX LowMemHiMemEMM FalseTrueOffOnNoYes LabelMovementFactor PointerSizePointerColorGrowth	ThresholdDelay SmallMediumLarge NormalReverseTransparent 	MouseTypeLanguageHorizontalSensitivityVerticalSensitivityDoubleThresholdActiveAccelerationProfileInterruptRateCursorDisplayDelayMemoryHardwareCursorSupportForceDefaultCursorRotationAnglePrimaryButtonSecondaryButton	ClickLock[AccelerationProfile1][AccelerationProfile2][AccelerationProfile3][AccelerationProfile4][DOSPointer][WindowsPointer]PhoenixBIOS BusSerialInportPS2MSX LowMemHiMemEMM FalseTrueOffOnNoYes LabelMovementFactor PointerSizePointerColorGrowth	ThresholdDelay SmallMediumLarge NormalReverseTransparent 	MouseTypeLanguageHorizontalSensitivityVerticalSensitivityDoubleThresholdActiveAccelerationProfileInterruptRateCursorDisplayDelayMemoryHardwareCursorSupportForceDefaultCursorRotationAnglePrimaryButtonSecondaryButton	ClickLock[AccelerationProfile1][AccelerationProfile2][AccelerationProfile3][AccelerationProfile4][DOSPointer][WindowsPointer]PhoenixBIOS BusSerialInportPS2MSX LowMemHiMemEMM FalseTrueOffOnNoYes LabelMovementFactor PointerSizePointerColorGrowth	ThresholdDelay SmallMediumLarge NormalReverseTransparent 	MouseTypeLanguageHorizontalSensitivityVerticalSensitivityDoubleThresholdActiveAccelerationProfileInterruptRateCursorDisplayDelayMemoryHardwareCursorSupportForceDefaultCursorRotationAnglePrimaryButtonSecondaryButton	ClickLock[AccelerationProfile1][AccelerationProfile2][AccelerationProfile3][AccelerationProfile4][DOSPointer][WindowsPointer]PhoenixBIOS BusSerialInportPS2MSX LowMemHiMemEMM FalseTrueOffOnNoYes LabelMovementFactor PointerSizePointerColorGrowth	ThresholdDelay SmallMediumLarge NormalReverseTransparent 	MouseTypeLanguageHorizontalSensitivityVerticalSensitivityDoubleThresholdActiveAccelerationProfileInterruptRateCursorDisplayDelayMemoryHardwareCursorSupportForceDefaultCursorRotationAnglePrimaryButtonSecondaryButton	ClickLock[AccelerationProfile1][AccelerationProfile2][AccelerationProfile3][AccelerationProfile4][DOSPointer][WindowsPointer]PhoenixBIOS BusSerialInportPS2MSX LowMemHiMemEMM FalseTrueOffOnNoYes LabelMovementFactor PointerSizePointerColorGrowth	ThresholdDelay SmallMediumLarge NormalReverseTransparent 	MouseTypeLanguageHorizontalSensitivityVerticalSensitivityDoubleThresholdActiveAccelerationProfileInterruptRateCursorDisplayDelayMemoryHardwareCursorSupportForceDefaultCursorRotationAnglePrimaryButtonSecondaryButton	ClickLock[AccelerationProfile1][AccelerationProfile2][AccelerationProfile3][AccelerationProfile4][DOSPointer][WindowsPointer]PhoenixBIOS BusSerialInportPS2MSX LowMemHiMemEMM FalseTrueOffOnNoYes LabelMovementFactor PointerSizePointerColorGrowth	ThresholdDelay SmallMediumLarge NormalReverseTransparent                                                                                                                                                                                                                                                                                        N��N�+ǋ�+�+�t���N����;L�v�L��6N�N��>L� t)L��ˋJ��ִ?�!r
����;>N�r��Ë߇�� rG<tC<
t?����3Ҋ�< t2��&�<Zw<Ar �$��Zw��Ar�� :�uGF�܋��Ë�����ɋ��Á�N�tN�<]tF�7 <=uF����;6N�s�<
t<u�;6N�s�<
t�<t�N�ÿN��6N���s��;6N�r��sì< t�<	t�N��SQ3��ǹ �� u��- ���, &�=�ǿ  ��Y�ً���� t� � �&�= u�[��[��3�&8t*V&�G< v�<;t�O&�< tG<;t
< v�FA��� ^����SVW���؎��� t�O&�G<\t&�\G��C< u�_^[��" r���� �6N��؎��D�Ëָ =�!ø >�!ËJ��B3ɋ��!r�� u�L��J�� B�!���PWV�N���rH��n�� �4�J�r��t���N����s��)��r$����n���4�$�r��=  t� �῁n����^_XÌ؎��r-�j�=  t%�J����N��B�r� ��s��J��P��� �3Zþ�n�� �4���r��r�� u�l� ��u��� ��w���u��u�n��u�4re���@�\��u�"rS�.Z�l�I��w��?��u�r5�C�/��w�$r(��À�u�7r�����u���u�� r�C� ���N������3ɬ<0r<9w,0��������r	Ȁ� r��$�<Ht<Ar<FvN;�Ë�3Ɋ�<0r�<9v$�<Ar�<Fw�,7�,0���������r����V���3Ҁ<.t��tJ�ѱ��<.u?F3ɬ<0r7<9w3,0��������ج<0r<9w,0ج<0r<9v�R�ñ��d 3���ZЋ�;�Ë���n���4�Q�r��Ë���n���4�>�r�� u�%Z ���u��t��� w�  ����u��%Z���u���tڃ�wո  ����u��%Z���u�%Z  �Ë���n���4���r�W���tl��u��dwc�)Z�Y���u��dwQ�*Z�Z���u��dw?�+Z�J���u��w-�� t(�-ZI�������u���,Z�
�t���/Z�M��@�t���u	�J�1Z���uI��w�Fي'�&E�I��w
�Fي�D��ʈ���߿��2����  ��  �2�� ���s�rU�N���rM��n��
�4���r,�@�r'�� u>�9��< t�� <t<
t<;t�����4�r뿻����I�:u�c �������� ����u)�|�t�
�u����? s��2������< t:O�v̈����t�
�u��I��? s��2�����< t:O�v����VW����< t6�����2������  ������|	�  �������	� ������_^��x�rH�N���r@����n���4���r)�C�r$�� u,�9 ����n���4���r�9�:�r���N����.��N�����u�: ����n���4��rԈ:����u�; �4�r��;���u�@ �Y�t��� t���dw��@��< �> �8�t΃� tɃ�dw���<�>�s��3n� ����)n���(�r�V���� s�ô0�!<rL.�, ��3�����I�� te&�= u��&�= tV���� �O��\�� ������+ο���������� �؎����C��!<w�A�E:�E\���)n�
 󤾠���� EnglishFrenchDutchGermanSwedishFinnishSpanish
PortugueseItalian �a��|���������� ������ܐ�$�8�T�ɒ�����'�X�l�������*�D�[�������1��L�^�x�����ԗ�e��������Ù���$������ƛ����(�<�X�͝�����+�\�p������.�H�_�����	MouseTypeLanguageHorizontalSensitivityVerticalSensitivityDoubleThresholdActiveAccelerationProfileInterruptRateCursorDisplayDelayMemoryHardwareCursorSupportForceDefaultCursorRotationAnglePrimaryButtonSecondaryButton	ClickLock[AccelerationProfile1][AccelerationProfile2][AccelerationProfile3][AccelerationProfile4][DOSPointer][WindowsPointer]PhoenixBIOS BusSerialInportPS2MSX LowMemHiMemEMM FalseTrueOffOnNoYes LabelMovementFactor PointerSizePointerColorGrowth	ThresholdDelay SmallMediumLarge NormalReverseTransparent 	MouseTypeLanguageHorizontalSensitivityVerticalSensitivityDoubleThresholdActiveAccelerationProfileInterruptRateCursorDisplayDelayMemoryHardwareCursorSupportForceDefaultCursorRotationAnglePrimaryButtonSecondaryButton	ClickLock[AccelerationProfile1][AccelerationProfile2][AccelerationProfile3][AccelerationProfile4][DOSPointer][WindowsPointer]PhoenixBIOS BusSerialInportPS2MSX LowMemHiMemEMM FalseTrueOffOnNoYes LabelMovementFactor PointerSizePointerColorGrowth	ThresholdDelay SmallMediumLarge NormalReverseTransparent 	MouseTypeLanguageHorizontalSensitivityVerticalSensitivityDoubleThresholdActiveAccelerationProfileInterruptRateCursorDisplayDelayMemoryHardwareCursorSupportForceDefaultCursorRotationAnglePrimaryButtonSecondaryButton	ClickLock[AccelerationProfile1][AccelerationProfile2][AccelerationProfile3][AccelerationProfile4][DOSPointer][WindowsPointer]PhoenixBIOS BusSerialInportPS2MSX LowMemHiMemEMM FalseTrueOffOnNoYes LabelMovementFactor PointerSizePointerColorGrowth	ThresholdDelay SmallMediumLarge NormalReverseTransparent 	MouseTypeLanguageHorizontalSensitivityVerticalSensitivityDoubleThresholdActiveAccelerationProfileInterruptRateCursorDisplayDelayMemoryHardwareCursorSupportForceDefaultCursorRotationAnglePrimaryButtonSecondaryButton	ClickLock[AccelerationProfile1][AccelerationProfile2][AccelerationProfile3][AccelerationProfile4][DOSPointer][WindowsPointer]PhoenixBIOS BusSerialInportPS2MSX LowMemHiMemEMM FalseTrueOffOnNoYes LabelMovementFactor PointerSizePointerColorGrowth	ThresholdDelay SmallMediumLarge NormalReverseTransparent 	MouseTypeLanguageHorizontalSensitivityVerticalSensitivityDoubleThresholdActiveAccelerationProfileInterruptRateCursorDisplayDelayMemoryHardwareCursorSupportForceDefaultCursorRotationAnglePrimaryButtonSecondaryButton	ClickLock[AccelerationProfile1][AccelerationProfile2][AccelerationProfile3][AccelerationProfile4][DOSPointer][WindowsPointer]PhoenixBIOS BusSerialInportPS2MSX LowMemHiMemEMM FalseTrueOffOnNoYes LabelMovementFactor PointerSizePointerColorGrowth	ThresholdDelay SmallMediumLarge NormalReverseTransparent 	MouseTypeLanguageHorizontalSensitivityVerticalSensitivityDoubleThresholdActiveAccelerationProfileInterruptRateCursorDisplayDelayMemoryHardwareCursorSupportForceDefaultCursorRotationAnglePrimaryButtonSecondaryButton	ClickLock[AccelerationProfile1][AccelerationProfile2][AccelerationProfile3][AccelerationProfile4][DOSPointer][WindowsPointer]PhoenixBIOS BusSerialInportPS2MSX LowMemHiMemEMM FalseTrueOffOnNoYes LabelMovementFactor PointerSizePointerColorGrowth	ThresholdDelay SmallMediumLarge NormalReverseTransparent 	MouseTypeLanguageHorizontalSensitivityVerticalSensitivityDoubleThresholdActiveAccelerationProfileInterruptRateCursorDisplayDelayMemoryHardwareCursorSupportForceDefaultCursorRotationAnglePrimaryButtonSecondaryButton	ClickLock[AccelerationProfile1][AccelerationProfile2][AccelerationProfile3][AccelerationProfile4][DOSPointer][WindowsPointer]PhoenixBIOS BusSerialInportPS2MSX LowMemHiMemEMM FalseTrueOffOnNoYes LabelMovementFactor PointerSizePointerColorGrowth	ThresholdDelay SmallMediumLarge NormalReverseTransparent 	MouseTypeLanguageHorizontalSensitivityVerticalSensitivityDoubleThresholdActiveAccelerationProfileInterruptRateCursorDisplayDelayMemoryHardwareCursorSupportForceDefaultCursorRotationAnglePrimaryButtonSecondaryButton	ClickLock[AccelerationProfile1][AccelerationProfile2][AccelerationProfile3][AccelerationProfile4][DOSPointer][WindowsPointer]PhoenixBIOS BusSerialInportPS2MSX LowMemHiMemEMM FalseTrueOffOnNoYes LabelMovementFactor PointerSizePointerColorGrowth	ThresholdDelay SmallMediumLarge NormalReverseTransparent 	MouseTypeLanguageHorizontalSensitivityVerticalSensitivityDoubleThresholdActiveAccelerationProfileInterruptRateCursorDisplayDelayMemoryHardwareCursorSupportForceDefaultCursorRotationAnglePrimaryButtonSecondaryButton	ClickLock[AccelerationProfile1][AccelerationProfile2][AccelerationProfile3][AccelerationProfile4][DOSPointer][WindowsPointer]PhoenixBIOS BusSerialInportPS2MSX LowMemHiMemEMM FalseTrueOffOnNoYes LabelMovementFactor PointerSizePointerColorGrowth	ThresholdDelay SmallMediumLarge NormalReverseTransparent                                                                                                                                                                                                                                                                                        ���+ǋ�+�+�t�������;�v���6���>� t)��ˋ��ִ?�!r
����;>�r��Ë߇�� rG<tC<
t?����3Ҋ�< t2��&�<Zw<Ar �$��Zw��Ar�� :�uGF�܋��Ë�����ɋ��Á��tN�<]tF�7 <=uF����;6�s�<
t<u�;6�s�<
t�<t�N�ÿ��6���s��;6�r��sì< t�<	t�N��SQ3��ǹ �� u��- ���, &�=�ǿ  ��Y�ً���� t� � �&�= u�[��[��3�&8t*V&�G< v�<;t�O&�< tG<;t
< v�FA��� ^����SVW���؎��� t�O&�G<\t&�\G��C< u�_^[��" r���� �6��؎��D�Ëָ =�!ø >�!Ë��B3ɋ��!r�� u����� B�!���PWV����rH�J��� �4�J�r��t�������s��)��r$���J����4�$�r��=  t� ��J�����^_X� &,28?EKQX^[mouse]
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         ���������������������������������U����Ȏ؎��|�� 2���=  u	�s�}�����< u����$$�E$���3ɴ<�!rݣz�����! ���F�؋v����N
�~
r�N
�~
v�F
 ���ؿ���s� �J��� �4�"�r]�q�rX����|�;6�t�< t�N�ο�+ϋ�����>y� t���y� ��r'V�2^N�<]u�y�<=uJ;6�tD�<;t<0s��
���;6�t0��>y� u�;6�t!�<t<
u�>y� u�;6�t
�<t�<
t�N�� ru���0�r�M�3۾J��� �4���S�2䀿|� u!�r���N�<]t�=���V� ^�� ��[C;^
rȋz���������ִA�!�؎�������V�!]����r�r�r&�����3�&�����3ɴ<�!r!&���غp����ش@�	 �!� B��3ɋ��!ô@�z������+��!�2仒�ڊ�� u�J����4P$����X���< t���Ju�J����4����w����u�J����4�JtJtJu��C���w���u�J����4=  t� ���v� J��W�'���_��3�V�J���
�4�[^�=���� �C< t������ V�J���
�4�5^�=�� ���2� ��2��-C���� V�J���
�4�	^�=��⠊��2� ���LC���q���r,;6�w&�bW��V�J��� �4��s
�����r��^_��6�w��tJt� �1�*��+�V�J����4� ^�=��V�J����4� ^�� V�J����4�u ^�=��GV�J����4�b ^�� � V�J����4�O ^�=��GV��^�� � V�J����4�1 ^�=��G�6 � � V�J����4� ^�=��G� � ��u�n�Ë�����������Q='s=�s=d s=
 s&�-3ҹ'��0���3ҹ���0���3ҹd ��0��±
��0���0�Y�2�P�����������.�X$S�`�؊[��	w�0�G��댰��
�È��WV�F�؋v���������² �����  ��Ƅ �  ������ �^_�VP��s�����trF�<�t���<�u��X^ð �1�>-��F������ �>OwP���X������P������P2������������$��>N t	��%$��
����A �t�A�t�A �>E t��Ҩt���t���t�� � t��2���t@��t���P"
Ȉ3҈C�6<�>>�Ĩ t(�u���6 �>�C����6��>��C�t(�u�
�6�>�C���6�>�CY[8Nt������>-��FF�ְ����������$��ְ����������������
ŘP�ְ���ׄ����ф$��ְ���ń���迄����������
ŘP��3��C���Њ��A �t�A �t�A�>E t����t���t���6<�>>��������"��ѻP"
ц8t&w���6 �>�C����6��>��C���"��ѻP"
��8t&w�
�6�>�C���6�>�CY[�-��惊�����݃������u4�L
�t �@u2���H�LC:Ms#� �1����H�L�@u��H �L �݀>� u� �K$�>H��0
�P�B�>C tD��<t%�< u�E
D��$<��"�:�u���<u��
�t��$�< t
>E�D��"�X2�>A�>Et�� �>Dt���H$�
ĢH�#�H�&H�$0�A�Et�H �Dt�H�6<�>>�C �H���"��ѻP"
��8t&w���6 �>�C����6��>��C�H������"��ѻP"
��8t&w�
�6�>�C���6�>�C2��H��������
I���2���������
J��Ȁ>� t�>K�����������L ��~ u��D�F��F,�^*�N(�>� u�� 
�y
�y$� �2��D��D� ¢Q��D��D���B�>C ta��t.�< u �E
D�Ҁ�<�������"�:�u���<u��
�t��$�< t�E������
�D�����������"�Ċ������A�@t�ˀ 2�E�������t���D�������t��$0
��)���z�����0�A�>E t��$���t��t�V2��
��4 � t�͉T2��t�ωR�C �Ћ6<�>>�"��ѻP"
ц8t&w���6 �>�C����6��>��C�"��ѻP"
��8t&w�
�6�>�C���6�>�C�Q��D�F��D�F��·�r r����j r����` r��ێûi�Q r�·�G r���3ۈ>��9 r���1 r��>C t����u�>��·� r��>w u%� ·� r���D��Ds
��u��t��X��D�F�2����������������֊���F�����F�ˀ>Q t��R�T�Q ���Ѳ���C�i�����۳���ƴs�f��� ������A�łƵ���̠����_��񴧶���=���� �m�1ş�����?���W����*�!��ݸ4�f�Ͼ[�3°�g���h�ˡ�.Ϸ�s�Y�@�\�+�.�����	���^��Ï�����E���~������W���i�n�˻½#�����&ĵ��-�i�D���`�>�3�k���������Q����T���7�yɉ˂��ϩҊէل��η�D��z�I�����S��ɢ���8�����'ښ���+���C���y��²�7�x�$���Ί�C�<֞گ�G�9�q�ܼr�ǿ��%���cƝ�~���W��ЕӜ�Invalid parameter
$Param�tre invalide
$Ongeldige parameter
$Ung�ltiger Parameter
$Ogiltig parameter
$Virheellinen parametri
$Par�metro no v�lido
$Par�metro inv�lido
$Parametro non valido
$Driver not installed -- Internal Error 1
$Gestionnaire non install� -- erreur interne 1
$Besturingsprogramma niet ge�nstalleerd -- Interne fout 1
$Treiber nicht installiert -- Interner Fehler 1
$Drivrutinen ej installerad -- Internt fel 1
$Ohjainta ei ole asennettu -- sis�inen virhe 1
$Controlador no instalado -- Error interno 1
$Controlador nao instalado -- Erro interno 1
$Driver non installato -- Errore interno 1
$Driver not installed -- Microsoft Mouse not found
$Gestionnaire non install� -- Microsoft Mouse introuvable
$Besturingsprogramma niet ge�nstalleerd -- Microsoft Muis niet gevonden
$Treiber nicht installiert -- Microsoft Mouse nicht gefunden
$Drivrutinen ej installerad -- Musen kunde ej hittas
$Ohjainta ei ole asennettu -- hiirt� ei l�ydy
$Controlador no instalado -- El Mouse no se encuentra
$Controlador nao instalado -- Mouse nao encontrado
$Driver non installato -- Mouse non trovato
$Driver not installed -- interrupt jumper missing
$Gestionnaire non install� -- cavalier
d'interruption introuvable
$Besturingsprogramma niet ge�nstalleerd -- Onderbrekingsspringer niet
aanwezig
$Treiber nicht installiert -- Interrupt-Jumper
nicht gefunden
$Drivrutinen ej installerad -- avbrottsbygel finns inte
$Ohjainta ei ole asennettu -- keskeytyksen kytkin puuttuu
$Controlador no instalado -- El puente de interrupci�n no se encuentra 
$Controlador nao instalado -- conector de interrup�ao nao encontrado
$Driver non installato -- ponticello di interrupt mancante
$Driver not installed -- multiple interrupt jumpers found
$Gestionnaire non install� -- plusieurs cavaliers
d'interruption pr�sents
$Besturingsprogramma niet ge�nstalleerd -- Meerdere
onderbrekingsspringers gevonden
$Treiber nicht installiert -- Mehrere Interrupt-Jumper gefunden
$Drivrutinen ej installerad -- multipla avbrottsbyglar
$Ohjainta ei ole asennettu -- liian monta keskeytyksen kytkint�
$Controlador no instalado -- Encontrados varios puentes de interrupci�n
$Controlador nao instalado -- m�ltiplos conectores de interrup�ao encontrados
$Driver non installato -- esiste pi� di un ponticello di interrupt
$MSX Mouse driver installed
$Le gestionnaire MSX Mouse est install�
$Microsoft MSX Mouse besturingsprogramma wordt ge�nstalleerd
$Maustreiber MSX installiert
$Drivrutinen installeras Microsoft MSX Mouse
$Asennetaan Microsoft MSX Mouse laiteohjain
$Controlador MSX del Mouse instalado
$Controlador do Microsoft MSX Mouse instalado
$Driver del MSX Mouse installato
$Mouse driver installed
$Gestionnaire de souris install�
$Microsoft Mouse besturingsprogramma wordt ge�nstalleerd
$Maustreiber installiert
$Installerar drivrutiner f�r Microsoft Mouse
$Asennetaan Microsoft Mouse laiteohjain
$Controlador del Mouse instalado
$Controlador do Microsoft Mouse instalado
$Driver del Microsoft Mouse installato
$Switch values passed to existing Mouse driver
$Param�tres transmis au gestionnaire existant de la souris
$Schakelwaarden doorgegeven naar bestaand besturingsprogramma
$Optionswerte an vorhandenen Maustreiber weitergeleitet
$Parameterv�rden flyttade till existerande drivrutin f�r musen
$Kytkinasetukset siirretty olemassaolevaan ohjaimeen
$Par�metros transferidos al controlador en uso
$Defini�oes passadas para o controlador existente do Mouse
$Parametri trasferiti al driver esistente
$Existing Mouse driver enabled
$Le gestionnaire existant de la souris est activ�
$Bestaand besturingsprogramma geactiveerd
$Vorhandener Maustreiber aktiviert
$Existerande drivrutin f�r musen aktiverad
$Olemassaoleva ohjain otetaan k�ytt��n
$El controlador en uso est� activado
$Controlador existente do Mouse ativado
$Driver esistente attivato
$Existing Mouse driver removed from memory
$Le gestionnaire existant de la souris est supprim� de la m�moire
$Bestaand besturingsprogramma uit geheugen verwijderd
$Vorhandener Maustreiber ist aus dem Speicher entfernt worden
$Existerande drivrutin avl�gsnad fr�n minnet
$Olemassaoleva ohjain poistettu muistista
$El controlador en uso fu� retirado de la memoria
$Controlador existente do Mouse retirado da mem�ria
$Driver esistente rimosso dalla memoria
$Existing Mouse driver disabled
$Le gestionnaire existant de la souris est d�sactiv�
$Bestaand besturingsprogramma inactief
$Vorhandener Maustreiber deaktiviert
$Existerande drivrutin inaktiverad
$Olemassaoleva ohjain poistetaan k�yt�st�
$El controlador del Mouse en uso est� desactivado
$Controlador existente do Mouse desativado
$Driver esistente disattivato
$Mouse Driver not installed
$Le gestionnaire de la souris n'est pas install�
$Besturingsprogramma niet ge�nstalleerd
$Maustreiber nicht installiert
$Drivrutinen ej installerad
$Ohjainta ei ole asennettu
$Controlador del Mouse no instalado
$Controlador do Mouse nao instalado
$Driver non installato
$Mouse driver installed, cannot change port (/i, /z, /c, and /b invalid)
$Le gestionnaire de la souris est install�, impossible de changer de
port (/i, /z, /c et /b invalides)
$Besturingsprogramma ge�nstalleerd, verandering van poort niet mogelijk
(/i, /z, /c en /b ongeldig)
$Maustreiber installiert, Anschlu� kann nicht gewechselt werden
(/i, /z, /c und /b ung�ltig)
$Drivrutinen installerad, kan inte byta port
(/i, /z, /c och /b ogiltiga)
$Ohjain asennettu, porttia ei voi vaihtaa
(virheellinen /i, /z, /c ja /b)
$Controlador del Mouse instalado,
no se puede cambiar el puerto (/i, /z, /c y /b no v�lidos)
$Controlador do Mouse instalado, nao � poss�vel mudar porta
(/i, /z, /c e /b inv�lidos)
$Driver installato, impossibile cambiare porta
(/i, /z, /c e /b non valide)
$Mouse driver already installed
$Le gestionnaire de la souris est d�j� install�
$Besturingsprogramma al ge�nstalleerd
$Maustreiber ist schon installiert
$Drivrutinen redan installerad
$Ohjain on jo asennettu
$Controlador del Mouse ya instalado
$Controlador do Mouse j� instalado
$Driver gi� installato
$Unable to disable Mouse driver -- Control Panel is active
$Impossible de d�sactiver le gestionnaire de la souris -- le Panneau
de configuration est actif
$Niet mogelijk besturingsprogramma uit te schakelen -- Configuratiescherm is
geactiveerd
$Maustreiber kann nicht deaktiviert werden -- Steuerungsfeld ist aktiv
$Kan inte inaktivera drivrutinen -- Kontrollpanelen �r aktiv
$Ohjainta ei voi poistaa k�yt�st� -- ohjaintaulu on aktiivinen
$No se puede desactivar el controlador -- El Panel de control est� activo
$Imposs�vel desativar controlador do Mouse -- painel de controle ativado
$Impossibile disattivare il driver -- Pannello di controllo in funzione
$Unable to disable Mouse driver -- Mouse Menu is active
$Impossible de d�sactiver le gestionnaire de la souris --
le menu souris est actif
$Niet mogelijk besturingsprogramma uit te schakelen -- Muismenu is geactiveerd
$Maustreiber kann nicht deaktiviert werden -- Mausmen� ist aktiv
$Kan inte inaktivera drivrutinen -- Musmenyn �r aktiv
$Ohjainta ei voi poistaa k�yt�st� -- hiirivalikko on aktiivinen
$No se puede desactivar el controlador del Mouse-- Un Men� del Mouse est� activo
$Imposs�vel desativar controlador do Mouse -- Menu do Mouse ativado
$Impossibile disattivare il driver -- Menu del Mouse in funzione
$Mouse driver installed.  Parameters /U, /E, /X no longer supported.
$Le gestionnaire de la souris est install�.
Les param�tres /U, /E, /X ne sont plus support�s.
$Muis besturingsprogramma ge�nstalleerd.
Parameters /U, /E en /X niet meer ondersteund.
$Maustreiber installiert. Parameter /U, /E, /X werden nicht mehr unterst�tzt.
$Drivrutinen installerad. Parametrar /U, /E, /X kan ej l�ngre anv�ndas.
$Hiiren ajuri asennettu.  Valitsimet /U, /E, /X ei en�� tuettu.
$Se ha instalado el controlador de Mouse.
No se aceptan m�s los par�metros /U, /E, /X.
$Controlador do Mouse instalado.  Os par�metros /U, /E, /X nao sao mais areitos.
$Driver installato.  Parametri /u, /e, /k non validi.
$Driver cannot be loaded from within Windows.  Exit Windows and try again.
$Le gestionnaire ne peut �tre charg� sous Windows.
Quittez Windows et essayez � nouveau.
$Besturingsprogramma kan niet vanuit Windows geladen worden.
Be�indig Windows en probeer opnieuw.
$Treiber kann nicht von Windows aus geladen werden.
Beenden Sie Windows und versuchen Sie es erneut.
$Drivrutinen kan ej laddas fr�n Windows.  Avsluta Windows och f�rs�k igen.
$Ajuria ei voi ladata Windowsista. Poistu Windowsista ja yrit� uudelleen.
$No se puede cargar el controlador desde Windows.
Salga de Windows y vuelva a intentar la operaci�n.
$O controlador nao pode ser carregado a partir do Windows.
Saia do Windows e tente novamente.
$Impossibile installare driver in una sessione di Windows.
Uscire Windows e riprovare.
$Microsoft (R) Mouse Driver Version 8.20
Copyright (C) Microsoft Corp. 1983-1992.  All rights reserved.
$Gestionnaire de la souris Microsoft (R) Mouse version 8.20
Copyright (C) Microsoft Corp. 1983-1992.  Tous droits r�serv�s.
$Microsoft (R) Mouse Besturingsprogramma Versie 8.20
Copyright (C) Microsoft Corp. 1983-1992.  Alle rechten voorbehouden.
$Microsoft (R) Mouse Treiber-Version 8.20
Copyright (C) 1983-1992 Microsoft Corp.  Alle Rechte vorbehalten.
$Microsoft (R) Mouse drivrutin version 8.20
(C) Copyright Microsoft Corporation 1983-1992. Med ensamr�tt.
$Microsoft (R) Mouse ohjainversio 8.20
(C) Copyright Microsoft Corporation 1983-1992. Kaikki oikeudet pid�tet��n.
$Controlador del Microsoft (R) Mouse Versi�n 8.20
Copyright Microsoft Corporation 1983-1992.  Todos los derechos reservados. 
$Controlador do Microsoft (R) Mouse Versao 8.20
Copyright (C) Microsoft Corp. 1983-1992.  Todos direitos reservados.
$Driver del Microsoft (R) Mouse Versione 8.20
Copyright (C) Microsoft Corp. 1983-1992.  Tutti i diritti sono riservati.
$Slow            Moderate        Fast            Unaccelerated   Faible          Moyenne         Maximale        Nulle           Langzaam        Gemiddeld       Snel            Onversneld      Niedrige        Mittlere        Hohe            Ohne            L�ngsam         Normal          Snabb           Oaccelererad    Hidas           Kohtuullinen    Nopea           Kiihdytt�m�t�n  Lento           Moderado        R�pido          No Acelerado    Devagar         Moderado        R�pido          Desacelerado    Lento           Medio           Veloce          Non accelerato  his problem.
;    Skip       Causes ScanDisk to skip fixing this problem, but continue
;               checking the disk.

   LostClust     = Prompt       ; Lost clusters
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        ;能够讲第二个扇区里面的内容加载到内存
;第一个程序mbr.asm,loader.asm


LOADER_BASE_ADDR equ 0x900 ;将loader放入0x900
LOADER_START_SECTOR equ 0x2 ;表示LBA方式,我们的loader存在第二块扇区

SECTION MBR vstart=0x7c00
	mov ax,cs   ;将代码段的地址0x7c00,放入计算寄存器
	mov ds,ax   ;将计算寄存器地址放入ds    ds=0x7c00  数据段寄存器
	mov es,ax	;将计算寄存器地址放入es    es=0x7c00  附加寄存器(额外寄存器)
	mov ss,ax	;将计算寄存器地址放入ss    ss=0x7c00  栈基址寄存器
	mov fs,ax	;将计算寄存器地址放入fs    fs=0x7c00  附加寄存器(额外寄存器)
	mov sp,0x7c00  ;将sp指向0x7c00
	mov ax,0xb800  ;ax指向显存的位置(文本模式的显示缓冲区)
	mov gs,ax   ;额外寄存器   将gs指向文本模式缓冲区

;调用10号中断
; AH = 0x06 功能
; AL = 0 表示全部清除
; BH = 上卷行的属性
; (CL,CH) 左上角 x,y
; (DL,DH) 右下角 x,y	
   mov ax,0600h  ;功能
   mov bx,0700h  ;通道号
   mov cx,0      ;左上角
   mov dx,184fh;(80,25)  文本模式就是80*25

   int 10h
;输入当前我们在MBR
   mov byte [gs:0x00],'1'
   mov byte [gs:0x01],0xA4

   mov byte [gs:0x02],' '
   mov byte [gs:0x03],0xA4

   mov byte [gs:0x04],'M'
   mov byte [gs:0x05],0xA4

   mov byte [gs:0x06],'B'
   mov byte [gs:0x07],0xA4

   mov byte [gs:0x08],'R'
   mov byte [gs:0x09],0xA4

   mov eax,LOADER_START_SECTOR   ;这是LBA读入的扇区
   mov bx,LOADER_BASE_ADDR       ;把mbr的基地址给起始寄存器
   mov cx,1                      ;要读取1个扇区
   call rd_disk                  ;读取扇区

   jmp LOADER_BASE_ADDR          ;跳到实际物理地址
rd_disk:
	;eax LBA的扇区号
	;bx  数据写入的内存地址
	;cx  读入的扇区数

	mov esi,eax   ;备份 eax  要读取的第2扇区
	mov di,cx   ;备份 cx     读取扇区数1
	;读写硬盘

	;设置读取的扇区数
	mov dx,0x1f2 ;读取第二个扇区
	mov al,cl    ;读取1个扇区
	out dx,al    ;把读取一个扇区放入dx

	mov eax,esi  ;恢复eax
	;将7-0位写入0x1f3
	mov dx,0x1f3
	out dx,al

	;将15-8位写给1f4
	mov cl,8
	shr eax,cl
	mov dx,0x1f4
	out dx,al

	;23-16位写给1f5
	shr eax,cl
	mov dx,0x1f5
	out dx,al

	;
	shr eax,cl
	and al,0x0f
	or al,0xe0  ;设置7-4位为1110,此时才是LBA模式
	mov dx,0x1f6
	out dx,al


	;向0x1f7写入读命令
	mov dx,0x1f7
	mov al,0x20
	out dx,al

	.not_ready:
	nop ;空指令
	in al,dx
	and al,0x88 ;硬盘准备好存储准备;7位为1表示硬盘忙

	cmp al,0x08 ;表示没准备好
	jnz .not_ready

	;读数据
	mov ax,di
	mov dx,256
	mul dx
	mov cx,ax
	mov dx,0x1f0

	.go_on:
		in ax,dx ;一个个读
		mov [bx],ax
		add bx,2
		loop .go_on
		ret

	times 510-($-$$) db 0	
	dw 0xaa55
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              conectix             ;� vpc   Wi2k    @      @  �?   ���raWo��ރP�ϓ$�                                                                                                                                                                                                                                                                                                                                                                                                                                            